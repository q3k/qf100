* NGSPICE file created from mkQF100Fabric.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__fakediode_2 abstract view
.subckt sky130_ef_sc_hd__fakediode_2 DIODE VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt mkQF100Fabric CLK RST_N cpu_ack_o cpu_adr_i[0] cpu_adr_i[10] cpu_adr_i[11]
+ cpu_adr_i[12] cpu_adr_i[13] cpu_adr_i[14] cpu_adr_i[15] cpu_adr_i[16] cpu_adr_i[17]
+ cpu_adr_i[18] cpu_adr_i[19] cpu_adr_i[1] cpu_adr_i[20] cpu_adr_i[21] cpu_adr_i[22]
+ cpu_adr_i[23] cpu_adr_i[24] cpu_adr_i[25] cpu_adr_i[26] cpu_adr_i[27] cpu_adr_i[28]
+ cpu_adr_i[29] cpu_adr_i[2] cpu_adr_i[30] cpu_adr_i[31] cpu_adr_i[3] cpu_adr_i[4]
+ cpu_adr_i[5] cpu_adr_i[6] cpu_adr_i[7] cpu_adr_i[8] cpu_adr_i[9] cpu_cyc_i cpu_dat_i[0]
+ cpu_dat_i[10] cpu_dat_i[11] cpu_dat_i[12] cpu_dat_i[13] cpu_dat_i[14] cpu_dat_i[15]
+ cpu_dat_i[16] cpu_dat_i[17] cpu_dat_i[18] cpu_dat_i[19] cpu_dat_i[1] cpu_dat_i[20]
+ cpu_dat_i[21] cpu_dat_i[22] cpu_dat_i[23] cpu_dat_i[24] cpu_dat_i[25] cpu_dat_i[26]
+ cpu_dat_i[27] cpu_dat_i[28] cpu_dat_i[29] cpu_dat_i[2] cpu_dat_i[30] cpu_dat_i[31]
+ cpu_dat_i[3] cpu_dat_i[4] cpu_dat_i[5] cpu_dat_i[6] cpu_dat_i[7] cpu_dat_i[8] cpu_dat_i[9]
+ cpu_dat_o[0] cpu_dat_o[10] cpu_dat_o[11] cpu_dat_o[12] cpu_dat_o[13] cpu_dat_o[14]
+ cpu_dat_o[15] cpu_dat_o[16] cpu_dat_o[17] cpu_dat_o[18] cpu_dat_o[19] cpu_dat_o[1]
+ cpu_dat_o[20] cpu_dat_o[21] cpu_dat_o[22] cpu_dat_o[23] cpu_dat_o[24] cpu_dat_o[25]
+ cpu_dat_o[26] cpu_dat_o[27] cpu_dat_o[28] cpu_dat_o[29] cpu_dat_o[2] cpu_dat_o[30]
+ cpu_dat_o[31] cpu_dat_o[3] cpu_dat_o[4] cpu_dat_o[5] cpu_dat_o[6] cpu_dat_o[7] cpu_dat_o[8]
+ cpu_dat_o[9] cpu_err_o cpu_rty_o cpu_sel_i[0] cpu_sel_i[1] cpu_sel_i[2] cpu_sel_i[3]
+ cpu_stb_i cpu_we_i gpio_ack_i gpio_adr_o[0] gpio_adr_o[10] gpio_adr_o[11] gpio_adr_o[12]
+ gpio_adr_o[13] gpio_adr_o[14] gpio_adr_o[15] gpio_adr_o[16] gpio_adr_o[17] gpio_adr_o[18]
+ gpio_adr_o[19] gpio_adr_o[1] gpio_adr_o[20] gpio_adr_o[21] gpio_adr_o[22] gpio_adr_o[23]
+ gpio_adr_o[24] gpio_adr_o[25] gpio_adr_o[26] gpio_adr_o[27] gpio_adr_o[28] gpio_adr_o[29]
+ gpio_adr_o[2] gpio_adr_o[30] gpio_adr_o[31] gpio_adr_o[3] gpio_adr_o[4] gpio_adr_o[5]
+ gpio_adr_o[6] gpio_adr_o[7] gpio_adr_o[8] gpio_adr_o[9] gpio_cyc_o gpio_dat_i[0]
+ gpio_dat_i[10] gpio_dat_i[11] gpio_dat_i[12] gpio_dat_i[13] gpio_dat_i[14] gpio_dat_i[15]
+ gpio_dat_i[16] gpio_dat_i[17] gpio_dat_i[18] gpio_dat_i[19] gpio_dat_i[1] gpio_dat_i[20]
+ gpio_dat_i[21] gpio_dat_i[22] gpio_dat_i[23] gpio_dat_i[24] gpio_dat_i[25] gpio_dat_i[26]
+ gpio_dat_i[27] gpio_dat_i[28] gpio_dat_i[29] gpio_dat_i[2] gpio_dat_i[30] gpio_dat_i[31]
+ gpio_dat_i[3] gpio_dat_i[4] gpio_dat_i[5] gpio_dat_i[6] gpio_dat_i[7] gpio_dat_i[8]
+ gpio_dat_i[9] gpio_dat_o[0] gpio_dat_o[10] gpio_dat_o[11] gpio_dat_o[12] gpio_dat_o[13]
+ gpio_dat_o[14] gpio_dat_o[15] gpio_dat_o[16] gpio_dat_o[17] gpio_dat_o[18] gpio_dat_o[19]
+ gpio_dat_o[1] gpio_dat_o[20] gpio_dat_o[21] gpio_dat_o[22] gpio_dat_o[23] gpio_dat_o[24]
+ gpio_dat_o[25] gpio_dat_o[26] gpio_dat_o[27] gpio_dat_o[28] gpio_dat_o[29] gpio_dat_o[2]
+ gpio_dat_o[30] gpio_dat_o[31] gpio_dat_o[3] gpio_dat_o[4] gpio_dat_o[5] gpio_dat_o[6]
+ gpio_dat_o[7] gpio_dat_o[8] gpio_dat_o[9] gpio_err_i gpio_rty_i gpio_sel_o[0] gpio_sel_o[1]
+ gpio_sel_o[2] gpio_sel_o[3] gpio_stb_o gpio_we_o ksc_ack_i ksc_adr_o[0] ksc_adr_o[10]
+ ksc_adr_o[11] ksc_adr_o[12] ksc_adr_o[13] ksc_adr_o[14] ksc_adr_o[15] ksc_adr_o[16]
+ ksc_adr_o[17] ksc_adr_o[18] ksc_adr_o[19] ksc_adr_o[1] ksc_adr_o[20] ksc_adr_o[21]
+ ksc_adr_o[22] ksc_adr_o[23] ksc_adr_o[24] ksc_adr_o[25] ksc_adr_o[26] ksc_adr_o[27]
+ ksc_adr_o[28] ksc_adr_o[29] ksc_adr_o[2] ksc_adr_o[30] ksc_adr_o[31] ksc_adr_o[3]
+ ksc_adr_o[4] ksc_adr_o[5] ksc_adr_o[6] ksc_adr_o[7] ksc_adr_o[8] ksc_adr_o[9] ksc_cyc_o
+ ksc_dat_i[0] ksc_dat_i[10] ksc_dat_i[11] ksc_dat_i[12] ksc_dat_i[13] ksc_dat_i[14]
+ ksc_dat_i[15] ksc_dat_i[16] ksc_dat_i[17] ksc_dat_i[18] ksc_dat_i[19] ksc_dat_i[1]
+ ksc_dat_i[20] ksc_dat_i[21] ksc_dat_i[22] ksc_dat_i[23] ksc_dat_i[24] ksc_dat_i[25]
+ ksc_dat_i[26] ksc_dat_i[27] ksc_dat_i[28] ksc_dat_i[29] ksc_dat_i[2] ksc_dat_i[30]
+ ksc_dat_i[31] ksc_dat_i[3] ksc_dat_i[4] ksc_dat_i[5] ksc_dat_i[6] ksc_dat_i[7] ksc_dat_i[8]
+ ksc_dat_i[9] ksc_dat_o[0] ksc_dat_o[10] ksc_dat_o[11] ksc_dat_o[12] ksc_dat_o[13]
+ ksc_dat_o[14] ksc_dat_o[15] ksc_dat_o[16] ksc_dat_o[17] ksc_dat_o[18] ksc_dat_o[19]
+ ksc_dat_o[1] ksc_dat_o[20] ksc_dat_o[21] ksc_dat_o[22] ksc_dat_o[23] ksc_dat_o[24]
+ ksc_dat_o[25] ksc_dat_o[26] ksc_dat_o[27] ksc_dat_o[28] ksc_dat_o[29] ksc_dat_o[2]
+ ksc_dat_o[30] ksc_dat_o[31] ksc_dat_o[3] ksc_dat_o[4] ksc_dat_o[5] ksc_dat_o[6]
+ ksc_dat_o[7] ksc_dat_o[8] ksc_dat_o[9] ksc_err_i ksc_rty_i ksc_sel_o[0] ksc_sel_o[1]
+ ksc_sel_o[2] ksc_sel_o[3] ksc_stb_o ksc_we_o spi_ack_i spi_adr_o[0] spi_adr_o[10]
+ spi_adr_o[11] spi_adr_o[12] spi_adr_o[13] spi_adr_o[14] spi_adr_o[15] spi_adr_o[16]
+ spi_adr_o[17] spi_adr_o[18] spi_adr_o[19] spi_adr_o[1] spi_adr_o[20] spi_adr_o[21]
+ spi_adr_o[22] spi_adr_o[23] spi_adr_o[24] spi_adr_o[25] spi_adr_o[26] spi_adr_o[27]
+ spi_adr_o[28] spi_adr_o[29] spi_adr_o[2] spi_adr_o[30] spi_adr_o[31] spi_adr_o[3]
+ spi_adr_o[4] spi_adr_o[5] spi_adr_o[6] spi_adr_o[7] spi_adr_o[8] spi_adr_o[9] spi_cyc_o
+ spi_dat_i[0] spi_dat_i[10] spi_dat_i[11] spi_dat_i[12] spi_dat_i[13] spi_dat_i[14]
+ spi_dat_i[15] spi_dat_i[16] spi_dat_i[17] spi_dat_i[18] spi_dat_i[19] spi_dat_i[1]
+ spi_dat_i[20] spi_dat_i[21] spi_dat_i[22] spi_dat_i[23] spi_dat_i[24] spi_dat_i[25]
+ spi_dat_i[26] spi_dat_i[27] spi_dat_i[28] spi_dat_i[29] spi_dat_i[2] spi_dat_i[30]
+ spi_dat_i[31] spi_dat_i[3] spi_dat_i[4] spi_dat_i[5] spi_dat_i[6] spi_dat_i[7] spi_dat_i[8]
+ spi_dat_i[9] spi_dat_o[0] spi_dat_o[10] spi_dat_o[11] spi_dat_o[12] spi_dat_o[13]
+ spi_dat_o[14] spi_dat_o[15] spi_dat_o[16] spi_dat_o[17] spi_dat_o[18] spi_dat_o[19]
+ spi_dat_o[1] spi_dat_o[20] spi_dat_o[21] spi_dat_o[22] spi_dat_o[23] spi_dat_o[24]
+ spi_dat_o[25] spi_dat_o[26] spi_dat_o[27] spi_dat_o[28] spi_dat_o[29] spi_dat_o[2]
+ spi_dat_o[30] spi_dat_o[31] spi_dat_o[3] spi_dat_o[4] spi_dat_o[5] spi_dat_o[6]
+ spi_dat_o[7] spi_dat_o[8] spi_dat_o[9] spi_err_i spi_rty_i spi_sel_o[0] spi_sel_o[1]
+ spi_sel_o[2] spi_sel_o[3] spi_stb_o spi_we_o vccd1 vssd1
XANTENNA__3140__A1 _5401_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4935__A _4935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3155_ _5719_/Q input43/X _3168_/S vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__mux2_2
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3691__A2 _4968_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _4316_/A _5392_/Q _3230_/S vssd1 vssd1 vccd1 vccd1 _4473_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4654__B _4654_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3050__S _3102_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4640__A1 _5464_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4670__A _4778_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _5068_/A vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _5737_/CLK _5727_/D vssd1 vssd1 vccd1 vccd1 _5727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2902__B _2902_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2939_ _2886_/Y _3455_/A _2938_/Y vssd1 vssd1 vccd1 vccd1 _3549_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__3286__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5658_ _5659_/CLK _5658_/D vssd1 vssd1 vccd1 vccd1 _5658_/Q sky130_fd_sc_hd__dfxtp_1
X_4609_ _4609_/A vssd1 vssd1 vccd1 vccd1 _5447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5589_ _5589_/CLK _5589_/D vssd1 vssd1 vccd1 vccd1 _5589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2706__A1 _2700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5651__D _5651_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3225__S _3235_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4548__C _4569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5006__A _5006_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3131__A1 input39/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5503__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input127_A ksc_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A1 _3756_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4283__C _4283_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__B2 _3851_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5653__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__B1 _2641_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4580__A _4580_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input92_A gpio_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3198__A1 _5341_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3196__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2945__A1 input2/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3627__C _4969_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output179_A _3746_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4739__B _4739_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3643__B _4988_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output346_A _3571_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5561__D _5561_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4458__C _4542_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3122__A1 _5398_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4177__D _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4755__A _4755_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4870__A1 _4101_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3673__A2 _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4870__B2 _4857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4960_ _4960_/A vssd1 vssd1 vccd1 vccd1 _5616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3911_ _3824_/X _3825_/X _3826_/X _3910_/Y vssd1 vssd1 vccd1 vccd1 _3911_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4891_ _4891_/A vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__buf_8
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4490__A _4595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3842_ _5772_/Q _3804_/X _3812_/X _3841_/Y vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__o22ai_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5736__D _5736_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3773_ _3763_/X _3766_/X _3768_/X _3772_/X _3331_/A vssd1 vssd1 vccd1 vccd1 _3773_/Y
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__2936__A1 _4431_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3820__B_N _3818_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5694_/CLK _5512_/D vssd1 vssd1 vccd1 vccd1 _5512_/Q sky130_fd_sc_hd__dfxtp_1
X_2724_ _2724_/A _2724_/B _2724_/C _2724_/D vssd1 vssd1 vccd1 vccd1 _2724_/Y sky130_fd_sc_hd__nand4_2
XFILLER_101_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5443_ _5531_/CLK _5443_/D vssd1 vssd1 vccd1 vccd1 _5443_/Q sky130_fd_sc_hd__dfxtp_1
X_2655_ _5377_/Q _2611_/A _2654_/Y vssd1 vssd1 vccd1 vccd1 _2782_/B sky130_fd_sc_hd__o21ai_4
Xoutput401 _3195_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput412 _3082_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__3834__A _4099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput423 _2892_/X vssd1 vssd1 vccd1 vccd1 spi_we_o sky130_fd_sc_hd__buf_2
X_5374_ _5765_/CLK _5374_/D vssd1 vssd1 vccd1 vccd1 _5374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2586_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2696_/A sky130_fd_sc_hd__buf_2
XANTENNA__4649__B _4649_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5526__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4325_ _4325_/A vssd1 vssd1 vccd1 vccd1 _5326_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5471__D _5471_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _5586_/Q vssd1 vssd1 vccd1 vccd1 _4256_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3113__A1 input36/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2884__S _3047_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3207_ _5728_/Q input53/X _3228_/S vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4665__A _4837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4187_ _4185_/X _4186_/Y _4846_/A vssd1 vssd1 vccd1 vccd1 _4187_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5676__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3138_ _5716_/Q input40/X _3186_/S vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2872__B1 _2544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3069_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3069_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4613__A1 _5450_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4613__B2 _4590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2913__A _3345_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5646__D _5646_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5381__D _5381_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4278__C _4278_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3104__A1 _5395_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4575__A _5204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3655__A2 _2927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4852__A1 _4836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__A2 _4074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3919__A _4110_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__C _4741_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__D _5556_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output296_A _3512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2918__A1 _2877_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3357__C _4697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5549__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2969__S _3246_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4469__B _4473_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3373__B _3380_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3894__A2 _3890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3092__C _4475_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4110_/A vssd1 vssd1 vccd1 vccd1 _4228_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5699__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__clkbuf_2
X_4041_ _4109_/A _4041_/B _4143_/C _4172_/D vssd1 vssd1 vccd1 vccd1 _4041_/X sky130_fd_sc_hd__and4_4
XANTENNA__4485__A _4485_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3820__C _3820_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4943_ _5156_/A vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4932__B _4940_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3829__A _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4874_ _4132_/X _4133_/X _4872_/X _4873_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _5577_/D
+ sky130_fd_sc_hd__o221a_1
X_3825_ _3857_/A vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5466__D _5466_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3756_ _3857_/A vssd1 vssd1 vccd1 vccd1 _3756_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2707_ _2707_/A vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__clkbuf_4
X_3687_ _4287_/A vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__buf_8
X_5426_ _5731_/CLK _5426_/D vssd1 vssd1 vccd1 vccd1 _5426_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput220 _3302_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[18] sky130_fd_sc_hd__buf_2
X_2638_ _2632_/Y _2613_/X _2932_/B vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__o21a_1
Xoutput231 _3324_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[28] sky130_fd_sc_hd__buf_2
Xoutput242 _3282_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput253 _3402_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[18] sky130_fd_sc_hd__buf_2
XANTENNA__3334__A1 _5491_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput264 _3437_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[28] sky130_fd_sc_hd__buf_2
X_5357_ _5737_/CLK _5357_/D vssd1 vssd1 vccd1 vccd1 _5357_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput275 _3370_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[9] sky130_fd_sc_hd__buf_2
X_2569_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput286 _3492_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput297 _3514_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[23] sky130_fd_sc_hd__buf_2
X_4308_ _4322_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__and2_1
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5288_ _5288_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5780_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3098__A0 _4320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4395__A _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4239_ _3806_/X _5689_/Q _4238_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2908__A _2908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4834__A1 _3733_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4834__B2 _4833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5003__B _5130_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3739__A _3757_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3270__B1 _4771_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4561__C _4569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5376__D _5376_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3177__C _4512_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3573__A1 _5605_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4289__B _4567_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input55_A cpu_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3876__A2 _3857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3089__A0 _5708_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2818__A _5377_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3640__C _4980_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output211_A _3256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output309_A _3474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5250__A1 _2665_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A2 _3804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3261__A0 _4386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__C _4485_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3800__A2 _3722_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5371__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3610_ _3613_/A _3620_/B _4957_/A vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__and3_1
XANTENNA__3087__C _4473_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4590_ _4590_/A vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3564__A1 _5603_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3995__B1_N _5465_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3541_ _3541_/A vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3384__A _3393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3472_ _3469_/X _3470_/X _4999_/C vssd1 vssd1 vccd1 vccd1 _3472_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5305__A2 _5268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5211_ _5211_/A vssd1 vssd1 vccd1 vccd1 _5735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3867__A2 _3848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5142_ _5142_/A vssd1 vssd1 vccd1 vccd1 _5706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5073_ _5666_/Q _4988_/A _3750_/X _5073_/B2 _5111_/B vssd1 vssd1 vccd1 vccd1 _5666_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2728__A _2728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4816__A1 _5548_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4816__B2 _4804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4024_ _3989_/X _5675_/Q _4023_/Y _3991_/X vssd1 vssd1 vccd1 vccd1 _4026_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2827__B1 _2658_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4943__A _5156_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__A1 _2592_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3559__A _3559_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5714__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4926_ _4938_/A _4938_/B _4926_/C vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__or3_1
XANTENNA__3252__A0 _4301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4857_ _5087_/A vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3808_ _4141_/A vssd1 vssd1 vccd1 vccd1 _3808_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4788_ _4788_/A vssd1 vssd1 vccd1 vccd1 _5533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2910__B _2910_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3739_ _3757_/A vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__buf_2
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3294__A _3316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _5446_/CLK _5409_/D vssd1 vssd1 vccd1 vccd1 _5409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3233__S _3233_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5014__A _5021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4556__C _4569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5394__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3469__A _3530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4035__A2 _3915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__A0 _5124_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3546__A1 _5598_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3408__S _3435_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output259_A _3421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3932__A _4139_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4747__B _4756_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2548__A _2652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3143__S _3168_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4274__A2 _3690_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4185__D _4185_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5737__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4763__A _4771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3234__A0 _5205_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5760_ _5766_/CLK _5760_/D vssd1 vssd1 vccd1 vccd1 _5760_/Q sky130_fd_sc_hd__dfxtp_1
X_2972_ _2876_/X _2882_/X _4552_/A vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4711_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4731_/B sky130_fd_sc_hd__buf_2
XANTENNA__2588__A2 _2574_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3785__A1 _5089_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5694_/CLK _5691_/D vssd1 vssd1 vccd1 vccd1 _5691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4642_ _4651_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _5465_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4573_ _4592_/A _5431_/Q _4665_/D _4573_/D vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__and4_1
XANTENNA__5744__D _5744_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2745__C1 _2574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3524_ _3526_/A _5656_/Q vssd1 vssd1 vccd1 vccd1 _3525_/A sky130_fd_sc_hd__and2_1
XANTENNA__4003__A _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4938__A _4938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3455_ _3455_/A vssd1 vssd1 vccd1 vccd1 _4289_/D sky130_fd_sc_hd__buf_6
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3386_ _4335_/B _5505_/Q _3400_/S vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3053__S _3248_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5056_ _5056_/A _5659_/Q _5056_/C _5056_/D vssd1 vssd1 vccd1 vccd1 _5057_/A sky130_fd_sc_hd__and4_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _4153_/A vssd1 vssd1 vccd1 vccd1 _4007_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3473__A0 _4392_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4673__A _4743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4392__B _4392_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4017__A2 _3848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3289__A _3289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3225__A0 _4368_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3776__A1 _3751_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4909_ _4913_/A _4913_/B _4909_/C vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__or3_1
XFILLER_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2921__A _5058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5654__D _5654_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3228__S _3228_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5009__A _5033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4848__A _4848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input157_A spi_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3902__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4583__A _4583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A cpu_adr_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3464__B1 _4995_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4661__C1 _4621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4008__A2 _4642_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2831__A _2831_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3646__B _4988_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2990__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__D _5564_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output376_A _3041_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3138__S _3186_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4192__A1 _3824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3365__C _4701_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2977__S _3252_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2742__A2 _2617_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4758__A _4771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3240_ _4292_/B _5383_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__mux2_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3171_ _3183_/A _3194_/B _4510_/C vssd1 vssd1 vccd1 vccd1 _3172_/A sky130_fd_sc_hd__and3_1
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3812__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4247__A2 _4660_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4493__A _4678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4924__C _4940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5739__D _5739_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3207__A0 _5728_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4404__C1 _4379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5743_ _5767_/CLK _5743_/D vssd1 vssd1 vccd1 vccd1 _5743_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4940__B _4940_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2955_ _5736_/Q input13/X _3228_/S vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__mux2_2
XFILLER_91_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2741__A _2741_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5674_ _5692_/CLK _5674_/D vssd1 vssd1 vccd1 vccd1 _5674_/Q sky130_fd_sc_hd__dfxtp_1
X_2886_ _2946_/A _5208_/A _2885_/X vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__o21ai_4
X_4625_ _5454_/Q _4623_/X _3782_/X _4660_/A vssd1 vssd1 vccd1 vccd1 _5454_/D sky130_fd_sc_hd__a211o_1
XFILLER_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5474__D _5474_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3048__S _5234_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4556_ _4556_/A _4556_/B _4569_/A vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__and3_1
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3507_ _3515_/A _5648_/Q vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__and2_1
XANTENNA__2733__A2 _4415_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4668__A _4668_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4487_ _4487_/A _4498_/B _4487_/C vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__or3_1
XANTENNA__3572__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3438_ _4368_/A _5520_/Q _3444_/S vssd1 vssd1 vccd1 vccd1 _4754_/C sky130_fd_sc_hd__mux2_1
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3376_/A _3380_/B _4705_/C vssd1 vssd1 vccd1 vccd1 _3370_/A sky130_fd_sc_hd__and3_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5108_ _5096_/X _4837_/A _4872_/A _5097_/X _4226_/B vssd1 vssd1 vccd1 vccd1 _5688_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5039_ _5043_/A _5649_/Q _5039_/C _5043_/D vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__and4_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2916__A _2916_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4643__C1 _4632_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5649__D _5649_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3749__A1 _2859_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3747__A _4091_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2651__A _2651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5432__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2972__A2 _2882_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5384__D _5384_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3921__A1 _3921_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4578__A _4600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5582__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3482__A _3482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4297__B _4310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput120 ksc_dat_i[1] vssd1 vssd1 vccd1 vccd1 _5065_/B2 sky130_fd_sc_hd__buf_2
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput131 ksc_dat_i[2] vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4882__C1 _4877_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput142 ksc_rty_i vssd1 vssd1 vccd1 vccd1 _3697_/B sky130_fd_sc_hd__clkbuf_1
Xinput153 spi_dat_i[18] vssd1 vssd1 vccd1 vccd1 _4097_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput164 spi_dat_i[28] vssd1 vssd1 vccd1 vccd1 _4242_/A1 sky130_fd_sc_hd__buf_2
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput175 spi_dat_i[9] vssd1 vssd1 vccd1 vccd1 _3937_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4229__A2 _4489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4744__C _4744_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5202__A _5202_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5559__D _5559_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3717__B1_N _5453_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4401__A2 _4400_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _2780_/A _2779_/A _2779_/C _2780_/D vssd1 vssd1 vccd1 vccd1 _2741_/B sky130_fd_sc_hd__nand4_2
XANTENNA__2561__A _5452_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3376__B _3380_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2671_ input20/X _2695_/B _2695_/C _2695_/D vssd1 vssd1 vccd1 vccd1 _2671_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4410_ _5228_/A vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__buf_8
XANTENNA__4165__A1 _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4165__B2 _4164_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5390_ _5435_/CLK _5390_/D vssd1 vssd1 vccd1 vccd1 _5390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _4341_/A vssd1 vssd1 vccd1 vccd1 _5333_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3912__A1 _3813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4488__A _4488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4272_ _3824_/X _3825_/X _3826_/X _4271_/Y vssd1 vssd1 vccd1 vccd1 _4272_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3223_ _5731_/Q input56/X _3223_/S vssd1 vssd1 vccd1 vccd1 _5200_/C sky130_fd_sc_hd__mux2_2
XFILLER_95_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3676__B1 _5589_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3154_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3183_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3428__A0 _4362_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2736__A _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3085_ _5143_/C _5322_/Q _3132_/S vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__mux2_8
XANTENNA__4625__C1 _4660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5469__D _5469_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4640__A2 _4639_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4951__A _4963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5455__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _4036_/A _5288_/A vssd1 vssd1 vccd1 vccd1 _3987_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3567__A _3622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3600__A0 _4344_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2938_ _2929_/Y _2937_/Y _5627_/Q vssd1 vssd1 vccd1 vccd1 _2938_/Y sky130_fd_sc_hd__o21ai_1
X_5726_ _5737_/CLK _5726_/D vssd1 vssd1 vccd1 vccd1 _5726_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2902__C _2902_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3286__B _5535_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5657_ _5659_/CLK _5657_/D vssd1 vssd1 vccd1 vccd1 _5657_/Q sky130_fd_sc_hd__dfxtp_1
X_2869_ _2859_/Y _3455_/A _5058_/B vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__a21oi_4
XFILLER_30_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4608_ _4611_/A _5447_/Q _5017_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__and4_1
X_5588_ _5694_/CLK _5588_/D vssd1 vssd1 vccd1 vccd1 _5588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2706__A2 _5266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4539_ _4539_/A vssd1 vssd1 vccd1 vccd1 _5418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3667__B1 _2845_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4864__C1 _4861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3419__A0 _4355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5022__A _5022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5379__D _5379_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A2 _4667_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4283__D _4283_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2642__A1 _2639_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4861__A _5268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5041__C1 _5023_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input85_A gpio_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4739__C _4739_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3643__C _4982_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3772__B_N _3770_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5328__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output241_A _3280_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3658__B1 _2845_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output339_A _3647_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3940__A _4147_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4870__A2 _4102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2556__A _5768_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3151__S _3151_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5478__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__A _4771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3968__A1_N _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3910_ _3905_/Y _3906_/X _3909_/Y vssd1 vssd1 vccd1 vccd1 _3910_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2633__A1 _2607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4890_ _5089_/A vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4278__B_N _3861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3841_ _3813_/X _3822_/Y _3839_/Y _3840_/X vssd1 vssd1 vccd1 vccd1 _3841_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_92_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3387__A _3393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3772_ _3769_/X _3770_/X _3772_/C _4278_/D vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__and4bb_1
X_5511_ _5555_/CLK _5511_/D vssd1 vssd1 vccd1 vccd1 _5511_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2936__A2 _4431_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2723_ _4439_/A _4439_/B _2782_/D _2787_/A _2787_/B vssd1 vssd1 vccd1 vccd1 _2724_/D
+ sky130_fd_sc_hd__o2111a_1
X_5442_ _5531_/CLK _5442_/D vssd1 vssd1 vccd1 vccd1 _5442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2654_ _2819_/A _2615_/X _2653_/Y _2736_/A vssd1 vssd1 vccd1 vccd1 _2654_/Y sky130_fd_sc_hd__o211ai_4
Xoutput402 _3201_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput413 _3088_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5373_ _5695_/CLK _5373_/D vssd1 vssd1 vccd1 vccd1 _5373_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5752__D _5752_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2585_ _2585_/A _2848_/B _2848_/C _2848_/D vssd1 vssd1 vccd1 vccd1 _2585_/Y sky130_fd_sc_hd__nand4_1
XFILLER_86_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4324_ _4324_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__or2_1
XFILLER_82_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4255_ _5482_/Q _4489_/A _4254_/X vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3649__B1 _4898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4946__A _4946_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3850__A _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__clkbuf_1
X_4186_ _2728_/A _3716_/X _5477_/Q vssd1 vssd1 vccd1 vccd1 _4186_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__4665__B _4665_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3137_ _3250_/S vssd1 vssd1 vccd1 vccd1 _3186_/S sky130_fd_sc_hd__buf_2
XANTENNA__3061__S _3230_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2872__A1 _5261_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3068_ _3092_/A _3073_/B _4464_/A vssd1 vssd1 vccd1 vccd1 _3069_/A sky130_fd_sc_hd__and3_1
XFILLER_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4613__A2 _4573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4681__A _4681_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3297__A _3303_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5709_ _5765_/CLK _5709_/D vssd1 vssd1 vccd1 vccd1 _5709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4129__A1 _4027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5662__D _5662_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5017__A _5021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4278__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4856__A _4872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__A _4115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5620__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4852__A2 _4837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__B1 _5573_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__C1 _4400_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5770__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3000__A _3000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2918__A2 _2879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output191_A _4137_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output289_A _3499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5572__D _5572_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3146__S _3146_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3879__B1 _3878_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4469__C _4469_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3373__C _4707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2985__S _3252_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4766__A _4766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4172_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4485__B _4500_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3820__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4056__B1 _4055_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__C1 _5238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4942_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5156_/A sky130_fd_sc_hd__buf_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4932__C _4940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5747__D _5747_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4873_ _5087_/A vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3824_ _3824_/A vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__buf_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__buf_4
XFILLER_101_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3845__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2706_ _2700_/X _5266_/A _2705_/Y vssd1 vssd1 vccd1 vccd1 _4439_/A sky130_fd_sc_hd__a21oi_1
X_3686_ _4196_/A vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__buf_4
X_5425_ _5435_/CLK _5425_/D vssd1 vssd1 vccd1 vccd1 _5425_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput210 _3949_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[9] sky130_fd_sc_hd__buf_2
X_2637_ _2637_/A _2637_/B _2637_/C vssd1 vssd1 vccd1 vccd1 _2932_/B sky130_fd_sc_hd__nand3_4
Xoutput221 _3304_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[19] sky130_fd_sc_hd__buf_2
XANTENNA__5482__D _5482_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput232 _3326_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[29] sky130_fd_sc_hd__buf_2
Xoutput243 _5805_/A vssd1 vssd1 vccd1 vccd1 gpio_cyc_o sky130_fd_sc_hd__buf_2
Xoutput254 _3406_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[19] sky130_fd_sc_hd__buf_2
X_5356_ _5737_/CLK _5356_/D vssd1 vssd1 vccd1 vccd1 _5356_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput265 _3440_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__5643__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2568_ _5382_/Q vssd1 vssd1 vccd1 vccd1 _2660_/A sky130_fd_sc_hd__inv_2
Xoutput276 _3448_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput287 _3494_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput298 _3516_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[24] sky130_fd_sc_hd__buf_2
X_4307_ _4307_/A vssd1 vssd1 vccd1 vccd1 _5318_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4676__A _4676_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5287_ _5287_/A vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4819__C1 _4805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4238_ _4238_/A vssd1 vssd1 vccd1 vccd1 _4238_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3098__A1 _5394_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2908__B _2908_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4834__A2 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5793__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4169_/A vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5003__C _5021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2924__A _3530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5300__A _5300_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3942__A_N _3832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3270__A1 _3267_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5657__D _5657_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3755__A _3755_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5392__D _5392_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4289__C _4407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input48_A cpu_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4586__A _5042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3490__A _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3089__A1 input63/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4286__B1 _4282_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2834__A _2902_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output204_A _3843_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__A _5223_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5250__A2 _2665_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3261__A1 _5526_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5567__D _5567_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5516__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4210__B1 _4200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3665__A _3665_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3540_ _3540_/A _3547_/B _4909_/C vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__and3_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5666__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3384__B _3397_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3471_ _4390_/A _5632_/Q _3645_/S vssd1 vssd1 vccd1 vccd1 _4999_/C sky130_fd_sc_hd__mux2_1
XFILLER_83_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5210_ _5223_/A _5215_/B _5210_/C vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__or3_1
XFILLER_83_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5141_ _5141_/A _5154_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__and3_1
XANTENNA__4496__A _4496_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _5072_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5665_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4816__A2 _4803_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _4023_/A vssd1 vssd1 vccd1 vccd1 _4023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2827__A1 _5759_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4029__B1 _4028_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5120__A _5120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5241__A2 _5227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4925_ _4925_/A vssd1 vssd1 vccd1 vccd1 _5601_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3252__A1 _5386_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5477__D _5477_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4856_ _4872_/A vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ _3807_/A vssd1 vssd1 vccd1 vccd1 _3807_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4787_ _4801_/A _5533_/Q _4796_/C vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__and3_1
XANTENNA__3575__A _3575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3738_ _4830_/B _3737_/X _5557_/Q vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2910__C _2910_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2763__B1 _2762_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__C1 _3959_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3669_ _4665_/B _3669_/B _4667_/A _4665_/C vssd1 vssd1 vccd1 vccd1 _3681_/B sky130_fd_sc_hd__nand4_4
XFILLER_66_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5408_ _5731_/CLK _5408_/D vssd1 vssd1 vccd1 vccd1 _5408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2919__A _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5339_ _5737_/CLK _5339_/D vssd1 vssd1 vccd1 vccd1 _5339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5014__B _5637_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5539__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input102_A gpio_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5387__D _5387_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__A1 _5314_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5689__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3485__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2754__B1 _2753_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2829__A _5369_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4747__C _4765_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5205__A _5223_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4259__B1 _4258_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output321_A _3592_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output419_A _3245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4763__B _4763_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2564__A _2622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _4388_/B _5423_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3234__A1 _5348_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ _4710_/A vssd1 vssd1 vccd1 vccd1 _5502_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A2 _3783_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5690_ _5690_/CLK _5690_/D vssd1 vssd1 vccd1 vccd1 _5690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ _4645_/A vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3395__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4572_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2745__B1 _2709_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3523_ _3523_/A vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3454_ _3281_/A _2899_/A _4679_/C vssd1 vssd1 vccd1 vccd1 _3454_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4938__B _4938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3385_ _3385_/A vssd1 vssd1 vccd1 vccd1 _3385_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5760__D _5760_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3334__S _3364_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3170__A0 _4346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5124_ _5128_/A _5143_/B _5124_/C vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__or3_1
XFILLER_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5658_/Q _5021_/D _3540_/A _5034_/A _5045_/X vssd1 vssd1 vccd1 vccd1 _5658_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4954__A _4954_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _3997_/X _3890_/X _4002_/X _4004_/X _4005_/X vssd1 vssd1 vccd1 vccd1 _4006_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_96_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3473__A1 _5633_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__C1 _2574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3225__A1 _5416_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _4908_/A vssd1 vssd1 vccd1 vccd1 _5595_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3776__A2 _5114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2984__A0 _5223_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4839_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__buf_6
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5670__D _5670_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3244__S _3252_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5025__A _5025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3161__A0 _5720_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5361__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3464__A1 _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4661__B1 _4254_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4413__B1 _4379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2975__A0 _5739_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2831__B _2831_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3419__S _3432_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3646__C _4984_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output271_A _3355_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4192__A2 _3857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output369_A _3028_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4758__B _4763_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4251__A2_N _5690_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2559__A _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5580__D _5580_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5704__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3170_ _4346_/A _5406_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _4510_/C sky130_fd_sc_hd__mux2_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4774__A _4774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4101__C1 _4100_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3207__A1 input53/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4404__B1 _2570_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5742_ _5766_/CLK _5742_/D vssd1 vssd1 vccd1 vccd1 _5742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2954_ _3250_/S vssd1 vssd1 vccd1 vccd1 _3228_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__4940__C _4940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2966__A0 _4386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5755__D _5755_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2741__B _2741_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5673_ _5697_/CLK _5673_/D vssd1 vssd1 vccd1 vccd1 _5673_/Q sky130_fd_sc_hd__dfxtp_1
X_2885_ _2700_/X _5266_/A _5349_/Q vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4624_ _4645_/A vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2718__B1 _2717_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4949__A _4949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4555_ _4555_/A vssd1 vssd1 vccd1 vccd1 _5424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3506_ _3517_/A vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__clkbuf_1
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _5397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5384__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3437_ _3437_/A vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5490__D _5490_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3143__A0 _5717_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3368_ _4324_/A _5500_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _4705_/C sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5099_/X _5094_/X _5066_/A _5102_/X _4214_/B vssd1 vssd1 vccd1 vccd1 _5687_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4684__A _4684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3299_ _3303_/A _5541_/Q vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__and2_1
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5038_ _5648_/Q _5033_/X _5029_/X _5034_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5648_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2916__B _2916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4643__B1 _4018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2654__C1 _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2932__A _2932_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3749__A2 _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5665__D _5665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3239__S _4375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4859__A _5081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5727__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__A _3763_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3921__A2 _4528_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3482__B _5637_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_10_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4189__A_N _3860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput110 ksc_dat_i[10] vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput121 ksc_dat_i[20] vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput132 ksc_dat_i[30] vssd1 vssd1 vccd1 vccd1 _4264_/B2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A cpu_adr_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4882__B1 _4207_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput143 spi_ack_i vssd1 vssd1 vccd1 vccd1 _3711_/A sky130_fd_sc_hd__buf_4
XFILLER_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput154 spi_dat_i[19] vssd1 vssd1 vccd1 vccd1 _4111_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput165 spi_dat_i[29] vssd1 vssd1 vccd1 vccd1 _4253_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput176 spi_err_i vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__buf_2
XFILLER_97_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5202__B _5202_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3003__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3938__A _4283_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2842__A _2842_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2948__A0 _5210_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5575__D _5575_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3149__S _3186_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3376__C _4709_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2670_ _5381_/Q _2691_/A _4441_/B vssd1 vssd1 vccd1 vccd1 _2779_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__2988__S _3229_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4165__A2 _4062_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4769__A _4769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4340_ _4344_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__and2_1
XANTENNA__3912__A2 _3904_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4271_ _4268_/Y _3828_/X _4270_/Y vssd1 vssd1 vccd1 vccd1 _4271_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3222_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3676__A1 _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3153_ _3153_/A vssd1 vssd1 vccd1 vccd1 _3153_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3612__S _3633_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3428__A1 _5517_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3084_ _3174_/A vssd1 vssd1 vccd1 vccd1 _3132_/S sky130_fd_sc_hd__buf_4
XANTENNA__2736__B _2736_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4625__B1 _3782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4951__B _4963_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3848__A _3848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3986_ _5780_/Q _3804_/X _3970_/X _3985_/Y vssd1 vssd1 vccd1 vccd1 _5288_/A sky130_fd_sc_hd__o22ai_4
XFILLER_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2939__B1 _2938_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5725_ _5737_/CLK _5725_/D vssd1 vssd1 vccd1 vccd1 _5725_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3600__A1 _5613_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2937_ _2937_/A _2937_/B _2937_/C _2937_/D vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__5485__D _5485_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3059__S _4375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2902__D _2902_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5656_ _5659_/CLK _5656_/D vssd1 vssd1 vccd1 vccd1 _5656_/Q sky130_fd_sc_hd__dfxtp_1
X_2868_ _3670_/A1 _2867_/X _5694_/Q vssd1 vssd1 vccd1 vccd1 _5058_/B sky130_fd_sc_hd__o21bai_4
X_4607_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5017_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4679__A _4699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5587_ _5589_/CLK _5587_/D vssd1 vssd1 vccd1 vccd1 _5587_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3364__A0 _4322_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4158__A2_N _5683_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2799_ _5590_/Q vssd1 vssd1 vccd1 vccd1 _2800_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4538_ _4538_/A _4550_/B _4538_/C vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__or3_1
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3116__A0 _4327_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4469_ _4487_/A _4473_/B _4469_/C vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__or3_1
XFILLER_28_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3667__A1 _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4864__B1 _4015_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2927__A _2927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3419__A1 _5514_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__A2 _2640_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3758__A _3758_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5041__B1 _5029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5395__D _5395_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4589__A _4600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input78_A gpio_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3493__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__C _3924_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3658__A1 _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output234_A _3328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3432__S _3432_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5213__A _5213_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3935__A2_N _5670_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output401_A _3195_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4771__B _4776_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2633__A2 _2617_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2572__A _5363_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _4153_/A vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__buf_4
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3387__B _3397_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3771_ _4099_/A vssd1 vssd1 vccd1 vccd1 _4278_/D sky130_fd_sc_hd__clkbuf_1
X_5510_ _5635_/CLK _5510_/D vssd1 vssd1 vccd1 vccd1 _5510_/Q sky130_fd_sc_hd__dfxtp_1
X_2722_ _5369_/Q _2565_/A _2721_/Y vssd1 vssd1 vccd1 vccd1 _2787_/B sky130_fd_sc_hd__o21ai_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5441_ _5446_/CLK _5441_/D vssd1 vssd1 vccd1 vccd1 _5441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4499__A _4499_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2653_ _2607_/X _2708_/A _5762_/Q vssd1 vssd1 vccd1 vccd1 _2653_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput403 _3206_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput414 _3093_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[6] sky130_fd_sc_hd__buf_2
X_2584_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2848_/D sky130_fd_sc_hd__clkbuf_4
X_5372_ _5695_/CLK _5372_/D vssd1 vssd1 vccd1 vccd1 _5372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4323_ _4323_/A vssd1 vssd1 vccd1 vccd1 _5325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4254_ _4254_/A _4265_/B _4254_/C vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__and3_1
XANTENNA__3649__A1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3205_ _3210_/A _3221_/B _4524_/C vssd1 vssd1 vccd1 vccd1 _3206_/A sky130_fd_sc_hd__and3_1
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2747__A _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3342__S _3364_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4185_ _4265_/A _4265_/B _4265_/C _4185_/D vssd1 vssd1 vccd1 vccd1 _4185_/X sky130_fd_sc_hd__and4_2
XANTENNA__5123__A _5223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4665__C _4665_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5422__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3136_ _3196_/A vssd1 vssd1 vccd1 vccd1 _3165_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2872__A2 _5261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3067_ _4308_/B _5389_/Q _3248_/S vssd1 vssd1 vccd1 vccd1 _4464_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4962__A _4962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4681__B _4681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__A _3578_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5572__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3297__B _5540_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ _4171_/A vssd1 vssd1 vccd1 vccd1 _4143_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5708_ _5766_/CLK _5708_/D vssd1 vssd1 vccd1 vccd1 _5708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4129__A2 _4095_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5639_ _5641_/CLK _5639_/D vssd1 vssd1 vccd1 vccd1 _5639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4202__A _4254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3888__A1 _3794_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5017__B _5639_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3252__S _3252_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5033__A _5033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4227__A_N _4075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input132_A ksc_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__A _4872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A1 _3961_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__B1 _4565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3488__A _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3576__A0 _4329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2918__A3 _2925_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output184_A _4036_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5208__A _5208_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4112__A _4145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3879__A1 _5458_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output351_A _5806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3951__A _3951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5445__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3162__S _3162_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4485__C _4485_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5595__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4782__A _4804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__B1 _4565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4056__B2 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4941_ _4941_/A vssd1 vssd1 vccd1 vccd1 _5609_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3398__A _3398_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4872_ _4872_/A vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3823_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _3823_/A vssd1 vssd1 vccd1 vccd1 _4628_/A sky130_fd_sc_hd__clkbuf_4
X_2705_ _5380_/Q vssd1 vssd1 vccd1 vccd1 _2705_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5763__D _5763_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3685_ _3685_/A _5270_/B _3685_/C vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__nand3_4
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5424_ _5731_/CLK _5424_/D vssd1 vssd1 vccd1 vccd1 _5424_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4022__A _4036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput200 _4263_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[29] sky130_fd_sc_hd__buf_2
X_2636_ input16/X _2761_/B _2647_/A _2761_/D vssd1 vssd1 vccd1 vccd1 _2637_/C sky130_fd_sc_hd__nand4b_2
Xoutput211 _3256_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput222 _3260_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput233 _3262_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput244 _3336_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4957__A _4957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5355_ _5737_/CLK _5355_/D vssd1 vssd1 vccd1 vccd1 _5355_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput255 _3340_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[1] sky130_fd_sc_hd__buf_2
X_2567_ _2707_/A _2549_/X _5746_/Q vssd1 vssd1 vccd1 vccd1 _2567_/Y sky130_fd_sc_hd__o21ai_1
Xoutput266 _3344_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__3861__A _4083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput277 _3450_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput288 _3497_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[15] sky130_fd_sc_hd__buf_2
X_4306_ _4306_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__or2_1
Xoutput299 _3519_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[25] sky130_fd_sc_hd__buf_2
XANTENNA__4676__B _4681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5286_ _5779_/Q _5269_/X _3953_/X _3964_/Y _5285_/X vssd1 vssd1 vccd1 vccd1 _5779_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4819__B1 _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4237_ _4263_/A _5306_/A vssd1 vssd1 vccd1 vccd1 _4237_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3072__S _3230_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2908__C _2908_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4168_ _4195_/A _4168_/B vssd1 vssd1 vccd1 vccd1 _4168_/Y sky130_fd_sc_hd__nor2_4
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4692__A _4692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3119_ _3179_/A vssd1 vssd1 vccd1 vccd1 _3168_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4099_ _4099_/A vssd1 vssd1 vccd1 vccd1 _4243_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5244__B1 _5751_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5300__B _5308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3270__A2 _3268_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5318__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3952__A1_N _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5673__D _5673_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3247__S _4375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5028__A _5028_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5468__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4289__D _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3771__A _4099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4286__A1 _5289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4286__B2 _4285_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2834__B _2908_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__B _5215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__A _4107_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3011__A _3011_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output399_A _3184_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3946__A _4153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4210__A1 _5794_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4210__B2 _4209_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2757__D1 _2806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3665__B _4128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5583__D _5583_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3384__C _4714_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3470_ _4295_/D vssd1 vssd1 vccd1 vccd1 _3470_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4777__A _4777_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3681__A _3742_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5140_ _5264_/C vssd1 vssd1 vccd1 vccd1 _5160_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4496__B _4500_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5069_/X _4890_/X _5070_/X _5045_/X _3812_/B vssd1 vssd1 vccd1 vccd1 _5664_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4022_ _4036_/A _5291_/A vssd1 vssd1 vccd1 vccd1 _4022_/Y sky130_fd_sc_hd__nor2_8
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2827__A2 _2683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4029__A1 _4029_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5758__D _5758_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5120__B _5130_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4924_ _4924_/A _4940_/B _4940_/C vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__and3_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4855_ _5090_/A vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2760__A _5361_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3806_ _3989_/A vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__buf_2
X_4786_ _4828_/A vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5610__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5493__D _5493_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3737_ _4003_/A vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__buf_2
XANTENNA__3067__S _3248_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2763__A1 _2760_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__B1 _3725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3668_ _2726_/A _3850_/A _5485_/Q vssd1 vssd1 vccd1 vccd1 _4665_/C sky130_fd_sc_hd__a21o_1
X_5407_ _5446_/CLK _5407_/D vssd1 vssd1 vccd1 vccd1 _5407_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4687__A _4687_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2619_ _2614_/Y _2615_/X _2618_/Y _2574_/A vssd1 vssd1 vccd1 vccd1 _2619_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_66_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5760__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3599_ _3599_/A vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3591__A _3594_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5338_ _5737_/CLK _5338_/D vssd1 vssd1 vccd1 vccd1 _5338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5269_ _5289_/A vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5014__C _5017_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2935__A _2935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5668__D _5668_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3766__A _3766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3485__B _5638_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2754__A1 _2569_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input60_A cpu_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4597__A _4597_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5205__B _5215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4259__A1 _4256_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3006__A _3006_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output314_A _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2845__A _5486_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4763__C _4763_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5221__A _5221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5578__D _5578_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2970_ _5217_/A _5353_/Q _3229_/S vssd1 vssd1 vccd1 vccd1 _4388_/B sky130_fd_sc_hd__mux2_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5633__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2580__A _2684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4640_ _5464_/Q _4639_/X _3973_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _5464_/D sky130_fd_sc_hd__a211o_1
XFILLER_89_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4571_ _5430_/Q _4563_/X _5807_/A _4564_/X _4565_/X vssd1 vssd1 vccd1 vccd1 _5430_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5783__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2745__A1 _5261_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3522_ _3526_/A _5655_/Q vssd1 vssd1 vccd1 vccd1 _3523_/A sky130_fd_sc_hd__and2_1
XFILLER_85_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3453_ _4301_/A _5490_/Q _3453_/S vssd1 vssd1 vccd1 vccd1 _4679_/C sky130_fd_sc_hd__mux2_1
XFILLER_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4938__C _4938_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2687__A_N _2734_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4300__A _4300_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3384_ _3393_/A _3397_/B _4714_/C vssd1 vssd1 vccd1 vccd1 _3385_/A sky130_fd_sc_hd__and3_1
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3170__A1 _5406_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5123_ _5223_/B vssd1 vssd1 vccd1 vccd1 _5143_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5054_ _5054_/A vssd1 vssd1 vccd1 vccd1 _5657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _4005_/A vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3350__S _3364_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5131__A _5131_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2681__B1 _2680_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5488__D _5488_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4970__A _4970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4907_ _4907_/A _4915_/B _4915_/C vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__and3_1
XFILLER_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3586__A _3622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2984__A1 _5356_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4838_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4769_ _4769_/A _4778_/B _4778_/C vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__and3_1
XFILLER_88_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5306__A _5306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3161__A1 input44/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5506__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2709__B1_N _5765_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2665__A _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3464__A2 _2927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4661__A1 _5482_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5656__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5398__D _5398_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4413__A1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3496__A _3504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2975__A1 input28/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2831__C _2848_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output264_A _3437_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3435__S _3435_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4758__C _4758_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5216__A _5216_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4215__B1_N _5479_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4101__B1 _3998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2575__A _5767_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3170__S _3204_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4790__A _4801_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4404__A1 _5361_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5741_ _5741_/CLK _5741_/D vssd1 vssd1 vccd1 vccd1 _5741_/Q sky130_fd_sc_hd__dfxtp_1
X_2953_ _3047_/A vssd1 vssd1 vccd1 vccd1 _3250_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2966__A1 _5422_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5672_ _5694_/CLK _5672_/D vssd1 vssd1 vccd1 vccd1 _5672_/Q sky130_fd_sc_hd__dfxtp_1
X_2884_ _5734_/Q input72/X _3047_/A vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__mux2_4
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4623_ _4652_/A vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2718__A1 _5368_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4554_ _4674_/A _4558_/B _4554_/C vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__or3_1
XFILLER_50_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4949__B _4965_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3505_ _3505_/A vssd1 vssd1 vccd1 vccd1 _3505_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5117__C1 _4848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5529__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4485_ _4485_/A _4500_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__and3_1
XANTENNA__5771__D _5771_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5126__A _5126_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3436_ _3445_/A _3445_/B _4751_/A vssd1 vssd1 vccd1 vccd1 _3437_/A sky130_fd_sc_hd__and3_1
XFILLER_63_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3143__A1 input41/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3407_/A vssd1 vssd1 vccd1 vccd1 _3396_/S sky130_fd_sc_hd__buf_2
XANTENNA__4965__A _4965_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5679__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5106_ _5096_/X _4837_/A _4872_/A _5097_/X _4200_/B vssd1 vssd1 vccd1 vccd1 _5686_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_100_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3298_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3298_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3080__S _3248_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4643__A1 _5466_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2916__C _2916_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2654__B1 _2653_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2932__B _2932_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2633__B1_N _5757_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2709__A1 _2616_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5108__C1 _4226_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5681__D _5681_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3255__S _3444_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__A3 _3714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5036__A _5043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input162_A spi_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput100 gpio_dat_i[4] vssd1 vssd1 vccd1 vccd1 _3862_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4875__A _5081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput111 ksc_dat_i[11] vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput122 ksc_dat_i[21] vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4882__A1 _4875_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput133 ksc_dat_i[31] vssd1 vssd1 vccd1 vccd1 _5112_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput144 spi_dat_i[0] vssd1 vssd1 vccd1 vccd1 _3718_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput155 spi_dat_i[1] vssd1 vssd1 vccd1 vccd1 _3782_/D sky130_fd_sc_hd__buf_2
Xinput166 spi_dat_i[2] vssd1 vssd1 vccd1 vccd1 _3796_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput177 spi_rty_i vssd1 vssd1 vccd1 vccd1 _3710_/A sky130_fd_sc_hd__buf_2
XANTENNA_input23_A cpu_adr_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5202__C _5208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3003__B _5433_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4398__B1 _4379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3938__B _4079_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2842__B _2842_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2948__A1 _5350_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3070__A0 _5705_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4115__A _4115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output381_A _2986_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3954__A _4128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4769__B _4778_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5591__D _5591_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_opt_3_1_CLK clkbuf_opt_3_1_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_1_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
X_4270_ _3829_/X _3830_/X _3831_/X _4269_/X _3836_/X vssd1 vssd1 vccd1 vccd1 _4270_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3221_ _3236_/A _3221_/B _4532_/A vssd1 vssd1 vccd1 vccd1 _3222_/A sky130_fd_sc_hd__and3_1
XANTENNA__3676__A2 _3736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3152_ _3152_/A _3165_/B _4500_/A vssd1 vssd1 vccd1 vccd1 _3153_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_9_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5531_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2884__A0 _5734_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _5707_/Q input62/X _3108_/S vssd1 vssd1 vccd1 vccd1 _5143_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4625__A1 _5454_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2736__C _2736_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4951__C _4951_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5766__D _5766_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3985_ _3813_/X _3974_/Y _3984_/Y _3946_/X vssd1 vssd1 vccd1 vccd1 _3985_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2939__A1 _2886_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3061__A0 _4306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5724_ _5737_/CLK _5724_/D vssd1 vssd1 vccd1 vccd1 _5724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2936_ _4431_/C _4431_/B _2821_/Y _2935_/Y vssd1 vssd1 vccd1 vccd1 _2937_/D sky130_fd_sc_hd__a211oi_4
XANTENNA__4025__A _4171_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4001__B_N _4000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5655_ _5659_/CLK _5655_/D vssd1 vssd1 vccd1 vccd1 _5655_/Q sky130_fd_sc_hd__dfxtp_1
X_2867_ _3697_/A _3697_/B vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__or2_2
XANTENNA__5351__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4606_ _5446_/Q _4589_/X _3062_/A _4590_/X _4598_/X vssd1 vssd1 vccd1 vccd1 _5446_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5586_ _5586_/CLK _5586_/D vssd1 vssd1 vccd1 vccd1 _5586_/Q sky130_fd_sc_hd__dfxtp_1
X_2798_ _3659_/A _3660_/A vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__or2_2
XANTENNA__4679__B _4688_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3364__A1 _5499_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _5417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4468_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__buf_2
XANTENNA__3116__A1 _5397_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4695__A _4695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3419_ _4355_/A _5514_/Q _3432_/S vssd1 vssd1 vccd1 vccd1 _4739_/C sky130_fd_sc_hd__mux2_2
XFILLER_28_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4399_ _5195_/A vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3667__A2 _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4864__A1 _4859_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2627__B1 _5743_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2943__A _3047_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__D _5676_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5041__A1 _5650_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5041__B2 _5034_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__B _5642_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3658__A2 _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5213__B _5225_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output227_A _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3014__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2618__B1 _5744_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3949__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2853__A _2853_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__C _4771_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5586__D _5586_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5374__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3387__C _4716_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3770_ _4000_/A vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ _2831_/A _2615_/X _2720_/Y _2699_/A _2672_/A vssd1 vssd1 vccd1 vccd1 _2721_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5440_ _5446_/CLK _5440_/D vssd1 vssd1 vccd1 vccd1 _5440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__buf_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput404 _3211_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[26] sky130_fd_sc_hd__buf_2
X_5371_ _5767_/CLK _5371_/D vssd1 vssd1 vccd1 vccd1 _5371_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput415 _3100_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[7] sky130_fd_sc_hd__buf_2
X_2583_ _2583_/A vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__buf_2
X_4322_ _4322_/A _4322_/B vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__and2_1
X_4253_ _4075_/A _4076_/A _4253_/C _4253_/D vssd1 vssd1 vccd1 vccd1 _4254_/C sky130_fd_sc_hd__and4bb_1
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3649__A2 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3623__S _3636_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3204_ _4360_/A _5412_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _4524_/C sky130_fd_sc_hd__mux2_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2857__B1 _5802_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4184_ _5685_/Q _4986_/A _3846_/X _4184_/B2 vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__a22oi_4
XANTENNA__2747__B _2779_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4665__D _4665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3135_ _3135_/A vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3066_ _5136_/A _5319_/Q _3102_/S vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__mux2_8
XANTENNA__5717__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3859__A _5561_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4681__C _4690_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5496__D _5496_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3968_ _3932_/X _5672_/Q _3967_/Y _3934_/X vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5765_/CLK _5707_/D vssd1 vssd1 vccd1 vccd1 _5707_/Q sky130_fd_sc_hd__dfxtp_1
X_2919_ _2919_/A vssd1 vssd1 vccd1 vccd1 _3699_/B sky130_fd_sc_hd__inv_2
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3594__A _3594_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3899_ _3806_/X _5668_/Q _3898_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _3900_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_30_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_24_CLK_A clkbuf_opt_2_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5638_ _5641_/CLK _5638_/D vssd1 vssd1 vccd1 vccd1 _5638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5569_ _5694_/CLK _5569_/D vssd1 vssd1 vccd1 vccd1 _5569_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4202__B _4228_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3888__A2 _3716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5017__C _5017_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5247__D1 _4429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A ksc_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5397__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__A1 _2709_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4065__A2 _4003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3769__A _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3273__A0 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input90_A gpio_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3576__A1 _5606_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5208__B _5225_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4112__B _4228_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3879__A2 _4444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3009__A _3009_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2848__A _2848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output344_A _3563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5224__A _5224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2839__B1 _5361_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4142__A2_N _5682_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5253__A1 _2657_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4940_ _4940_/A _4940_/B _4940_/C vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__and3_1
XANTENNA__2583__A _2583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4871_ _4859_/X _4860_/X _4119_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5576_/D sky130_fd_sc_hd__a211o_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3822_ _5456_/Q _3815_/X _3821_/X vssd1 vssd1 vccd1 vccd1 _3822_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_18_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _3848_/A vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ _2704_/A vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__buf_2
XANTENNA__4303__A _4441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3684_ _5801_/Q _3790_/A _4199_/A _5094_/A vssd1 vssd1 vccd1 vccd1 _3685_/C sky130_fd_sc_hd__nand4b_2
XFILLER_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5423_ _5435_/CLK _5423_/D vssd1 vssd1 vccd1 vccd1 _5423_/Q sky130_fd_sc_hd__dfxtp_1
X_2635_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2761_/D sky130_fd_sc_hd__clkbuf_4
Xoutput201 _3803_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4022__B _5291_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput212 _3285_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_86_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput223 _3307_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput234 _3328_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[30] sky130_fd_sc_hd__buf_2
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _5741_/CLK _5354_/D vssd1 vssd1 vccd1 vccd1 _5354_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput245 _3374_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2566_ input4/X vssd1 vssd1 vccd1 vccd1 _2761_/A sky130_fd_sc_hd__inv_4
Xoutput256 _3410_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__4957__B _4965_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput267 _3443_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _5317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput278 _3452_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[2] sky130_fd_sc_hd__buf_2
Xoutput289 _3499_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5285_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4819__A1 _5550_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3353__S _3441_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4819__B2 _4804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4676__C _4690_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5134__A _5134_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4236_ _5796_/Q _3747_/X _4226_/X _4235_/Y vssd1 vssd1 vccd1 vccd1 _5306_/A sky130_fd_sc_hd__o22ai_4
XFILLER_99_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2908__D _2908_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4973__A _5025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4167_ _5791_/Q _4091_/X _4159_/X _4166_/Y vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__o22ai_4
XFILLER_99_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5229__D1 _4377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3118_ _3118_/A vssd1 vssd1 vccd1 vccd1 _3118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _4098_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5244__A1 _2813_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3589__A _3589_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3255__A0 _4381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3049_ _3174_/A vssd1 vssd1 vccd1 vccd1 _3102_/S sky130_fd_sc_hd__buf_4
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3907__B_N _3833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5044__A _5044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4286__A2 _5800_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4883__A _5235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3499__A _3499_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3246__A0 _5700_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2834__C _2834_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__C _5210_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2850__B _2850_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output294_A _3508_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3438__S _3444_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4210__A2 _4070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2757__C1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5219__A _5223_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4123__A _4123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5412__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3681__B _3681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2578__A input6/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5562__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3173__S _3186_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4496__C _4512_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__buf_4
XFILLER_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4021_ _3747_/X _5782_/Q _4017_/Y _4020_/Y vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__4793__A _4801_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__A2 _3954_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4434__C1 _4310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5120__C _5236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4923_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4940_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4854_ _4836_/X _4837_/X _3944_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5566_/D sky130_fd_sc_hd__a211o_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3805_ _5068_/A vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__clkbuf_1
X_4785_ _3316_/A _4804_/A _3723_/X vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5774__D _5774_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5129__A _5129_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3736_ _3736_/A vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4217__A_N _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2763__A2 _2696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__A1 _3922_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4968__A _4968_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3667_ _2726_/A _3850_/A _2845_/X vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3872__A _5562_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5406_ _5731_/CLK _5406_/D vssd1 vssd1 vccd1 vccd1 _5406_/Q sky130_fd_sc_hd__dfxtp_1
X_2618_ _2616_/X _2617_/X _5744_/Q vssd1 vssd1 vccd1 vccd1 _2618_/Y sky130_fd_sc_hd__o21ai_2
X_3598_ _3613_/A _3601_/B _4951_/C vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__and3_1
XFILLER_66_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3591__B _3601_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5337_ _5731_/CLK _5337_/D vssd1 vssd1 vccd1 vccd1 _5337_/Q sky130_fd_sc_hd__dfxtp_1
X_2549_ _2549_/A vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__buf_2
XANTENNA__3083__S _3108_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5268_ _5268_/A _5268_/B _5268_/C _5268_/D vssd1 vssd1 vccd1 vccd1 _5768_/D sky130_fd_sc_hd__nor4_1
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4219_ _3735_/A _4003_/A _5583_/Q vssd1 vssd1 vccd1 vccd1 _4219_/X sky130_fd_sc_hd__o21a_2
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3476__B1 _5005_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5014__D _5021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5199_ _5199_/A vssd1 vssd1 vccd1 vccd1 _5730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2935__B _2935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3228__A0 _5732_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3112__A _3112_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5435__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5684__D _5684_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5039__A _5043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3400__A0 _4344_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2754__A2 _2544_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5585__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3782__A _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input53_A cpu_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5205__C _5205_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4259__A2 _4692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3467__A0 _4388_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5221__B _5225_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3219__A0 _5198_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output307_A _3468_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3022__A _3022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3957__A _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2861__A _5697_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5594__D _5594_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3168__S _3168_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _4570_/A vssd1 vssd1 vccd1 vccd1 _5429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ _3521_/A vssd1 vssd1 vccd1 vccd1 _3521_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2745__A2 _2615_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4788__A _4788_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3692__A _4138_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3452_ _3281_/A _2899_/A _4676_/A vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__o21a_1
XFILLER_100_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3383_ _4333_/A _5504_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _4714_/C sky130_fd_sc_hd__mux2_1
XFILLER_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5122_ _5195_/A vssd1 vssd1 vccd1 vccd1 _5223_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5056_/A _5657_/Q _5056_/C _5056_/D vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__and4_1
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3458__B1 _4990_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4655__C1 _4645_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4004_ _3961_/X _4003_/X _5569_/Q vssd1 vssd1 vccd1 vccd1 _4004_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5769__D _5769_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__A1 _2813_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5458__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5080__C1 _3936_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4906_ _4906_/A vssd1 vssd1 vccd1 vccd1 _5594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2771__A _2771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4837_ _4837_/A vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3078__S _3126_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4186__A1 _2728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4768_ _4768_/A vssd1 vssd1 vccd1 vccd1 _5526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4698__A _4698_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3719_ _3823_/A vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__clkbuf_4
X_4699_ _4699_/A _4714_/B _4699_/C vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__or3_1
XANTENNA__2631__A_N _2878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5306__B _5308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3107__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4894__C1 _4883_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3449__A0 _4297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2946__A _2946_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4646__C1 _4645_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2665__B _2665_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5679__D _5679_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4661__A2 _4652_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4413__A2 _2596_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3777__A _4057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5071__C1 _3812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3496__B _5643_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2831__D _2831_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3909__D1 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output257_A _3413_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3017__A _3017_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4885__C1 _4877_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3451__S _3451_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4637__C1 _4632_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5232__A _5232_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4101__A1 _4098_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5600__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5589__D _5589_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4790__B _5535_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4404__A2 _4400_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5062__C1 _3705_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3687__A _4287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5750__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2952_ _2876_/X _2882_/X _4545_/C vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3612__A0 _4351_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740_ _5766_/CLK _5740_/D vssd1 vssd1 vccd1 vccd1 _5740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2883_ _2544_/B _2708_/X _5266_/C vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__a21o_2
X_5671_ _5697_/CLK _5671_/D vssd1 vssd1 vccd1 vccd1 _5671_/Q sky130_fd_sc_hd__dfxtp_1
X_4622_ _4638_/A _4622_/B vssd1 vssd1 vccd1 vccd1 _5453_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2718__A2 _2613_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _5423_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3626__S _3633_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4949__C _4965_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3504_ _3504_/A _5647_/Q vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__and2_1
XANTENNA__4311__A _4311_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5117__B1 _5070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4484_ _4484_/A vssd1 vssd1 vccd1 vccd1 _5396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5126__B _5130_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3435_ _4366_/B _5519_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3679__B1 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3366_ _3366_/A vssd1 vssd1 vccd1 vccd1 _3366_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4965__B _4965_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5685_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3297_ _3303_/A _5540_/Q vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__and2_1
XFILLER_100_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5142__A _5142_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5036_ _5043_/A _5647_/Q _5039_/C _5043_/D vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__and4_1
XANTENNA__5499__D _5499_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4643__A2 _4639_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2916__D _2929_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4981__A _4981_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2654__A1 _2819_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2932__C _2932_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2709__A2 _2617_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5108__B1 _5097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5036__B _5647_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4867__C1 _4861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input155_A spi_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5623__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput101 gpio_dat_i[5] vssd1 vssd1 vccd1 vccd1 _3873_/C sky130_fd_sc_hd__clkbuf_2
Xinput112 ksc_dat_i[12] vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput123 ksc_dat_i[22] vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4882__A2 _4876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput134 ksc_dat_i[3] vssd1 vssd1 vccd1 vccd1 _3807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2676__A _2750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput145 spi_dat_i[10] vssd1 vssd1 vccd1 vccd1 _3956_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__3271__S _3451_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput156 spi_dat_i[20] vssd1 vssd1 vccd1 vccd1 _4130_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput167 spi_dat_i[30] vssd1 vssd1 vccd1 vccd1 _4265_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5292__C1 _5285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input16_A cpu_adr_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5773__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4891__A _4891_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3842__B1 _3812_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4398__A1 _2835_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3938__C _3938_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3300__A _3300_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2842__C _2842_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3070__A1 input60/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output374_A _3039_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4769__C _4778_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5227__A _5227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3970__A _4109_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4858__C1 _4843_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3220_ _4366_/B _5415_/Q _3230_/S vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3151_ _4340_/B _5403_/Q _3151_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2586__A _2621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2884__A1 input72/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3181__S _3192_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3082_ _3082_/A vssd1 vssd1 vccd1 vccd1 _3082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4086__B1 _4085_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5283__C1 _5310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4625__A2 _4623_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5035__C1 _5023_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4306__A _4306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3210__A _3210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3984_ _3940_/X _3825_/X _3975_/X _3983_/Y vssd1 vssd1 vccd1 vccd1 _3984_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2939__A2 _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5723_ _5737_/CLK _5723_/D vssd1 vssd1 vccd1 vccd1 _5723_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3061__A1 _5388_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2935_ _2935_/A _2935_/B _2935_/C vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__nand3_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5654_ _5659_/CLK _5654_/D vssd1 vssd1 vccd1 vccd1 _5654_/Q sky130_fd_sc_hd__dfxtp_1
X_2866_ _2877_/A _2879_/A _2866_/C _2866_/D vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__nand4_4
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _5445_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5782__D _5782_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3356__S _3364_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2797_ _2853_/B _2853_/C _2797_/C vssd1 vssd1 vccd1 vccd1 _3403_/A sky130_fd_sc_hd__nand3_4
X_5585_ _5694_/CLK _5585_/D vssd1 vssd1 vccd1 vccd1 _5585_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4679__C _4679_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5137__A _5137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4041__A _4109_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5646__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4536_ _4536_/A _4556_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__and3_1
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4976__A _4990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4467_ _5270_/A vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__buf_2
XFILLER_28_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4849__C1 _4848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3418_ _3418_/A vssd1 vssd1 vccd1 vccd1 _3433_/B sky130_fd_sc_hd__clkbuf_1
X_4398_ _2835_/Y _2837_/X _4379_/X vssd1 vssd1 vccd1 vccd1 _5358_/D sky130_fd_sc_hd__o21ai_1
XFILLER_28_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4864__A2 _4860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input8_A cpu_adr_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3349_ _3349_/A vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__clkbuf_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5796__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3091__S _3248_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _5640_/Q _5010_/X _5806_/A _5011_/X _4823_/X vssd1 vssd1 vccd1 vccd1 _5640_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2627__A1 _2593_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5041__A2 _5033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5692__D _5692_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5047__A _5056_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__A _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5213__C _5231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4068__B1 _4058_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3014__B _5438_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2618__A1 _2616_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3949__B _5284_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2853__B _2853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5519__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3030__A _3038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4100__A_N _3999_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _2593_/X _2594_/X _5754_/Q vssd1 vssd1 vccd1 vccd1 _2720_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5669__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3684__B _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2651_ _2651_/A vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__clkinv_4
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3176__S _3209_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2694__B1_N _5755_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput405 _3217_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[27] sky130_fd_sc_hd__buf_2
X_2582_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2848_/C sky130_fd_sc_hd__buf_4
X_5370_ _5800_/CLK _5370_/D vssd1 vssd1 vccd1 vccd1 _5370_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput416 _3106_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _4321_/A vssd1 vssd1 vccd1 vccd1 _5324_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4796__A _4801_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4252_ _4252_/A _4252_/B _4252_/C _4664_/A vssd1 vssd1 vccd1 vccd1 _4252_/X sky130_fd_sc_hd__and4_4
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3203_ _5191_/C _5342_/Q _3234_/S vssd1 vssd1 vccd1 vccd1 _4360_/A sky130_fd_sc_hd__mux2_8
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4195_/A _5302_/A vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__nor2_4
XFILLER_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2857__A1 _2560_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3205__A _3210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2747__C _2779_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3134_ _3152_/A _3134_/B _4494_/C vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__and3_1
XFILLER_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3065_ _5704_/Q input57/X _5234_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5777__D _5777_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4036__A _4036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _3967_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5706_ _5766_/CLK _5706_/D vssd1 vssd1 vccd1 vccd1 _5706_/Q sky130_fd_sc_hd__dfxtp_1
X_2918_ _2877_/A _2879_/A _2925_/C _5660_/Q vssd1 vssd1 vccd1 vccd1 _2919_/A sky130_fd_sc_hd__a31oi_4
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3898_ _3898_/A vssd1 vssd1 vccd1 vccd1 _3898_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3594__B _3601_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2793__B1 _2792_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5637_ _5641_/CLK _5637_/D vssd1 vssd1 vccd1 vccd1 _5637_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3086__S _3230_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2849_ _5745_/Q _2577_/X _2848_/Y _2565_/A vssd1 vssd1 vccd1 vccd1 _2850_/D sky130_fd_sc_hd__o211ai_2
XFILLER_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5568_ _5586_/CLK _5568_/D vssd1 vssd1 vccd1 vccd1 _5568_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4202__C _4202_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4519_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5017__D _5021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5499_ _5538_/CLK _5499_/D vssd1 vssd1 vccd1 vccd1 _5499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__C1 _4848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__A _3250_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__A2 _5261_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A ksc_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3273__A1 _5530_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5687__D _5687_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_2_1_CLK clkbuf_opt_2_1_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_1_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4222__B1 _4214_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input83_A gpio_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2784__B1 _2661_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5208__C _5208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4112__C _4112_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3733__C1 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2848__B _2848_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2839__A1 _2809_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output337_A _3545_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3025__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5341__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2864__A _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__A2 _2658_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5597__D _5597_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4870_ _4101_/X _4102_/X _4856_/X _4857_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _5575_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5491__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3821_ _4283_/A _4283_/B _3821_/C vssd1 vssd1 vccd1 vccd1 _3821_/X sky130_fd_sc_hd__and3_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4213__B1 _4212_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3695__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3752_ _4147_/A _4062_/A _3678_/X _3662_/Y vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__o22ai_1
XFILLER_18_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2703_ _4417_/C _4417_/B _2689_/Y _2702_/Y vssd1 vssd1 vccd1 vccd1 _2724_/C sky130_fd_sc_hd__a211oi_1
X_3683_ _3683_/A vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__buf_4
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5422_ _5731_/CLK _5422_/D vssd1 vssd1 vccd1 vccd1 _5422_/Q sky130_fd_sc_hd__dfxtp_1
X_2634_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2761_/B sky130_fd_sc_hd__clkbuf_4
Xoutput202 _4275_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput213 _3287_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput224 _3309_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[21] sky130_fd_sc_hd__buf_2
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput235 _3330_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[31] sky130_fd_sc_hd__buf_2
X_2565_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__clkbuf_4
X_5353_ _5737_/CLK _5353_/D vssd1 vssd1 vccd1 vccd1 _5353_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput246 _3377_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput257 _3413_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[21] sky130_fd_sc_hd__buf_2
XANTENNA__4957__C _4965_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput268 _3446_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[31] sky130_fd_sc_hd__buf_2
X_4304_ _4322_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__and2_1
Xoutput279 _3454_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_88_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _5284_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5778_/D sky130_fd_sc_hd__nand2_1
XANTENNA__4819__A2 _4803_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4235_ _3792_/D _4229_/Y _4234_/Y _4153_/X vssd1 vssd1 vccd1 vccd1 _4235_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_29_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4166_ _4059_/X _4654_/B _4165_/Y _3840_/X vssd1 vssd1 vccd1 vccd1 _4166_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__5229__C1 _5228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2774__A _4830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3117_ _3123_/A _3134_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__and3_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4097_ _4097_/A1 _3954_/X _3994_/X _4096_/Y vssd1 vssd1 vccd1 vccd1 _4649_/B sky130_fd_sc_hd__a31oi_4
XFILLER_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5150__A _5150_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5244__A2 _2831_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3048_ _5702_/Q input35/X _5234_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3255__A1 _5524_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4999_ _5128_/A _5005_/B _4999_/C vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__or3_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2766__B1 _2850_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2949__A _2949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3191__A0 _5725_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5364__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2684__A _2684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5060__A _5094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3246__A1 input69/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__B1 _4402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2834__D _2834_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2850__C _2850_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2757__B1 _2595_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5219__B _5223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4123__B _5297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output287_A _3494_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2859__A _5660_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5707__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3182__A0 _4351_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5235__A _5235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3681__C _3681_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _3707_/X _4019_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _4020_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4793__B _5537_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2594__A _2652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__A3 _3994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4434__B1 _4433_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4922_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4940_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ _3925_/X _3926_/X _4832_/X _4833_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _5565_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3629__S _3636_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3804_ _4070_/A vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__buf_4
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4314__A _4385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4784_ _5532_/Q _4780_/X _5805_/A _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _5532_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3945__C1 _3944_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3735_ _3735_/A vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__buf_2
XFILLER_31_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3960__A2 _3958_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5405_ _5446_/CLK _5405_/D vssd1 vssd1 vccd1 vccd1 _5405_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5387__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2617_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__buf_4
XANTENNA__5790__D _5790_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3364__S _3364_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3597_ _4342_/A _5612_/Q _3597_/S vssd1 vssd1 vccd1 vccd1 _4951_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3173__A0 _5722_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5145__A _5145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3591__C _4945_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5336_ _5737_/CLK _5336_/D vssd1 vssd1 vccd1 vccd1 _5336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2548_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__buf_4
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4984__A _4990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5267_ _5267_/A vssd1 vssd1 vccd1 vccd1 _5767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _4098_/X _3958_/A _4781_/A _4217_/X vssd1 vssd1 vccd1 vccd1 _4218_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3476__A1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5198_ _5198_/A _5202_/B _5208_/C vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__and3_1
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4149_ _4082_/X _4083_/X _4149_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _4149_/X sky130_fd_sc_hd__and4bb_1
XFILLER_84_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2935__C _2935_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3228__A1 input58/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2987__A0 _5742_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3539__S _3642_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4224__A _4224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2739__B1 _4421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5039__B _5649_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3400__A1 _5509_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2754__A3 _2549_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3782__B _4283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2679__A _2679_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3164__A0 _4344_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input46_A cpu_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3467__A1 _5631_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3303__A _3303_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5221__C _5231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3219__A1 _5345_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output202_A _4275_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2978__B1 _4554_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3449__S _3453_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3927__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3973__A _4145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3520_ _3526_/A _5654_/Q vssd1 vssd1 vccd1 vccd1 _3521_/A sky130_fd_sc_hd__and2_1
XFILLER_89_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3451_ _4299_/B _5489_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2589__A _2794_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3155__A0 _5719_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3382_ _3418_/A vssd1 vssd1 vccd1 vccd1 _3397_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _5121_/A vssd1 vssd1 vccd1 vccd1 _5698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4104__C1 _4007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5052_ _5656_/Q _5021_/D _3540_/A _5034_/A _5045_/X vssd1 vssd1 vccd1 vccd1 _5656_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3458__A1 _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4655__B1 _4174_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4003_/A vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4309__A _4309_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3863__D1 _3836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__A2 _2615_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2969__A0 _5738_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5080__B1 _5076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4905_ _4913_/A _4913_/B _4905_/C vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__or3_1
XFILLER_55_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5785__D _5785_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4044__A _4145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4836_ _5081_/A vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4186__A2 _3716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4979__A _4979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4767_ _4771_/A _4776_/B _4767_/C vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__or3_1
XANTENNA__3883__A _3883_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4591__C1 _4576_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3718_ _3718_/A1 _4528_/A _3714_/X _3717_/Y vssd1 vssd1 vccd1 vccd1 _4622_/B sky130_fd_sc_hd__a31oi_4
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4698_ _4698_/A vssd1 vssd1 vccd1 vccd1 _5497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3649_ _3469_/X _3470_/X _4898_/A vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3146__A0 _4338_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4894__B1 _4872_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5319_ _5766_/CLK _5319_/D vssd1 vssd1 vccd1 vccd1 _5319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3449__A1 _5488_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4646__B1 _4044_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2665__C _2665_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5402__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5071__B1 _5045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input100_A gpio_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5695__D _5695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3269__S _3444_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5552__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3909__C1 _3907_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4889__A _5081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3793__A _3849_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4885__B1 _4233_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4637__B1 _3938_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4101__A2 _3958_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output417_A _3112_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3033__A _3033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4790__C _4796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5062__B1 _5061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2951_ _4381_/A _5420_/Q _3235_/S vssd1 vssd1 vccd1 vccd1 _4545_/C sky130_fd_sc_hd__mux2_1
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3612__A1 _5616_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4270__D1 _3836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5670_ _5694_/CLK _5670_/D vssd1 vssd1 vccd1 vccd1 _5670_/Q sky130_fd_sc_hd__dfxtp_1
X_2882_ _2882_/A vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2820__C1 _2606_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__clkbuf_2
X_4552_ _4552_/A _4556_/B _4569_/A vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__and3_1
XFILLER_89_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3503_ _3503_/A vssd1 vssd1 vccd1 vccd1 _3503_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5117__A1 _5696_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5117__B2 _4847_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4483_ _4487_/A _4498_/B _4483_/C vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__or3_1
XANTENNA__3128__A0 _4331_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3434_ _3434_/A vssd1 vssd1 vccd1 vccd1 _3434_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5126__C _5236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__A1 _3979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4030__C _4030_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3365_ _3376_/A _3380_/B _4701_/A vssd1 vssd1 vccd1 vccd1 _3366_/A sky130_fd_sc_hd__and3_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__S _3642_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4965__C _4965_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5425__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5104_ _5096_/X _5089_/X _5090_/X _5097_/X _4172_/B vssd1 vssd1 vccd1 vccd1 _5684_/D
+ sky130_fd_sc_hd__a311o_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3296_ _3296_/A vssd1 vssd1 vccd1 vccd1 _3296_/X sky130_fd_sc_hd__clkbuf_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5646_/Q _5033_/X _5029_/X _5034_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5646_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2654__A2 _2615_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5575__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__A _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2782__A _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3089__S _3126_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2932__D _2932_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4205__C _4205_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4819_ _5550_/Q _4803_/X _3339_/A _4804_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5550_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5799_ _5800_/CLK _5799_/D vssd1 vssd1 vccd1 vccd1 _5799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4502__A _4558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5108__A1 _5096_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3118__A _3118_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5036__C _5039_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4867__B1 _4050_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2957__A _3174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput102 gpio_dat_i[6] vssd1 vssd1 vccd1 vccd1 _3891_/C sky130_fd_sc_hd__buf_2
Xinput113 ksc_dat_i[13] vssd1 vssd1 vccd1 vccd1 _5086_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput124 ksc_dat_i[23] vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4126__A1_N _3989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput135 ksc_dat_i[4] vssd1 vssd1 vccd1 vccd1 _3847_/B2 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input148_A spi_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4619__B1 _4971_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput146 spi_dat_i[11] vssd1 vssd1 vccd1 vccd1 _3972_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput157 spi_dat_i[21] vssd1 vssd1 vccd1 vccd1 _4144_/C sky130_fd_sc_hd__clkbuf_1
Xinput168 spi_dat_i[31] vssd1 vssd1 vccd1 vccd1 _4283_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5292__B1 _4026_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3842__A1 _5772_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3788__A _3788_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3842__B2 _3841_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2692__A _5370_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4398__A2 _2837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4412__A _4412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output367_A _3024_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3028__A _3028_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5448__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__B1 _4856_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3970__B _3970_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2867__A _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3150_ _5169_/A _5333_/Q _3162_/S vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__mux2_8
XFILLER_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5598__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3081_ _3092_/A _3105_/B _4471_/A vssd1 vssd1 vccd1 vccd1 _3082_/A sky130_fd_sc_hd__and3_1
XFILLER_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4086__A1 _4081_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5283__B1 _3918_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3698__A _3698_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5035__B1 _5029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4306__B _4310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3983_ _3976_/Y _3906_/X _3982_/Y vssd1 vssd1 vccd1 vccd1 _3983_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3597__A0 _4342_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3210__B _3221_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5722_ _5741_/CLK _5722_/D vssd1 vssd1 vccd1 vccd1 _5722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2934_ _4439_/A _4439_/B _2782_/A _2779_/B _2779_/D vssd1 vssd1 vccd1 vccd1 _2937_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_17_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5653_ _5659_/CLK _5653_/D vssd1 vssd1 vccd1 vccd1 _5653_/Q sky130_fd_sc_hd__dfxtp_1
X_2865_ _2917_/A _2917_/B vssd1 vssd1 vccd1 vccd1 _2866_/D sky130_fd_sc_hd__nor2_1
X_4604_ _4611_/A _5445_/Q _4604_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__and4_1
XANTENNA__4322__A _4322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5584_ _5586_/CLK _5584_/D vssd1 vssd1 vccd1 vccd1 _5584_/Q sky130_fd_sc_hd__dfxtp_1
X_2796_ _2796_/A _2796_/B _2796_/C vssd1 vssd1 vccd1 vccd1 _2797_/C sky130_fd_sc_hd__nor3_2
XFILLER_89_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4535_ _4535_/A vssd1 vssd1 vccd1 vccd1 _5416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4041__B _4041_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4466_ _4466_/A vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__buf_8
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4976__B _4990_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4849__B1 _3864_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3417_ _3417_/A vssd1 vssd1 vccd1 vccd1 _3417_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2777__A _5556_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3372__S _3400_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4397_ _4397_/A vssd1 vssd1 vccd1 vccd1 _5357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5153__A _5153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3348_ _3357_/A _3361_/B _4688_/C vssd1 vssd1 vccd1 vccd1 _3349_/A sky130_fd_sc_hd__and3_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4992__A _4992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3279_ _3281_/A _5532_/Q vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__and2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5018_ _5018_/A vssd1 vssd1 vccd1 vccd1 _5639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2627__A2 _2594_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3401__A _3412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5047__B _5653_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5740__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4068__A1 _5785_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__B2 _4067_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2618__A2 _2617_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4407__A _4407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3311__A _3311_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2853__C _2853_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3030__B _5445_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3457__S _3645_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5238__A _5238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3684__C _4199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2650_ _2650_/A _2650_/B vssd1 vssd1 vccd1 vccd1 _2780_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2581_ _2581_/A vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__clkbuf_2
Xoutput406 _3222_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput417 _3112_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[9] sky130_fd_sc_hd__buf_2
X_4320_ _4320_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__or2_1
XANTENNA__3751__B1 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4796__B _5539_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2597__A _2622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4251_ _4139_/X _5690_/Q _4250_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _4252_/B sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__3192__S _3192_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3202_ _5727_/Q input52/X _3223_/S vssd1 vssd1 vccd1 vccd1 _5191_/C sky130_fd_sc_hd__mux2_2
X_4182_ _5792_/Q _4070_/X _4172_/X _4181_/Y vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__2857__A2 _2949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__B _3221_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2747__D _2782_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3133_ _4333_/A _5400_/Q _3146_/S vssd1 vssd1 vccd1 vccd1 _4494_/C sky130_fd_sc_hd__mux2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _4617_/A vssd1 vssd1 vccd1 vccd1 _3092_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4317__A _4317_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3221__A _3236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4036__B _4036_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3966_ _4036_/A _3966_/B vssd1 vssd1 vccd1 vccd1 _3966_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5613__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5705_ _5765_/CLK _5705_/D vssd1 vssd1 vccd1 vccd1 _5705_/Q sky130_fd_sc_hd__dfxtp_1
X_2917_ _2917_/A _2917_/B _2917_/C vssd1 vssd1 vccd1 vccd1 _2925_/C sky130_fd_sc_hd__nor3_4
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5793__D _5793_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3897_ _3949_/A _3897_/B vssd1 vssd1 vccd1 vccd1 _3897_/Y sky130_fd_sc_hd__nor2_8
XFILLER_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5148__A _5152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2793__A1 _5362_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5636_ _5641_/CLK _5636_/D vssd1 vssd1 vccd1 vccd1 _5636_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3594__C _4949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2848_ _2848_/A _2848_/B _2848_/C _2848_/D vssd1 vssd1 vccd1 vccd1 _2848_/Y sky130_fd_sc_hd__nand4_1
X_5567_ _5802_/CLK _5567_/D vssd1 vssd1 vccd1 vccd1 _5567_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4987__A _5056_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5763__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2779_ _2779_/A _2779_/B _2779_/C _2779_/D vssd1 vssd1 vccd1 vccd1 _2781_/A sky130_fd_sc_hd__nand4_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4518_ _4518_/A vssd1 vssd1 vccd1 vccd1 _5409_/D sky130_fd_sc_hd__clkbuf_1
X_5498_ _5538_/CLK _5498_/D vssd1 vssd1 vccd1 vccd1 _5498_/Q sky130_fd_sc_hd__dfxtp_1
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4558_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2702__D1 _2701_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__B1 _2716_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4222__A1 _5795_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4222__B2 _4221_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5058__A _5058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2784__A1 _2783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input76_A gpio_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4897__A _5025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5804__425 vssd1 vssd1 vccd1 vccd1 _5804__425/HI cpu_rty_o sky130_fd_sc_hd__conb_1
XFILLER_100_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3733__B1 _3725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_opt_2_1_CLK_A clkbuf_opt_2_1_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3306__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2848__C _2848_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5538_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2839__A2 _2750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3025__B _5443_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output232_A _3326_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2864__B _2864_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4137__A _4195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3041__A _3041_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5636__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3976__A _5568_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2880__A _2909_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3820_ _3817_/X _3818_/X _3820_/C _4043_/D vssd1 vssd1 vccd1 vccd1 _3821_/C sky130_fd_sc_hd__and4bb_1
XFILLER_18_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4213__B2 _3808_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3751_ _5662_/Q _5002_/A _3750_/X _5065_/B2 vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__5786__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3187__S _3219_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2702_ _2690_/Y _2903_/A _2932_/C _2932_/D _2701_/Y vssd1 vssd1 vccd1 vccd1 _2702_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3682_ _3682_/A vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__buf_4
X_5421_ _5435_/CLK _5421_/D vssd1 vssd1 vccd1 vccd1 _5421_/Q sky130_fd_sc_hd__dfxtp_1
X_2633_ _2607_/A _2617_/X _5757_/Q vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__o21bai_2
Xoutput203 _4287_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput214 _3289_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__4600__A _4600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5352_ _5737_/CLK _5352_/D vssd1 vssd1 vccd1 vccd1 _5352_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput225 _3311_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2564_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2565_/A sky130_fd_sc_hd__buf_4
Xoutput236 _3266_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput247 _3381_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput258 _3417_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[22] sky130_fd_sc_hd__buf_2
X_4303_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput269 _3349_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[3] sky130_fd_sc_hd__buf_2
X_5283_ _5777_/Q _5269_/X _3918_/X _3928_/Y _5310_/B vssd1 vssd1 vccd1 vccd1 _5777_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3216__A _3236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4234_ _4147_/X _3722_/X _3758_/A _4233_/Y vssd1 vssd1 vccd1 vccd1 _4234_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_96_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _3824_/A _4062_/X _4163_/X _4164_/X _4835_/A vssd1 vssd1 vccd1 vccd1 _4165_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__S _3654_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5229__B1 _2628_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _4327_/B _5397_/Q _3151_/S vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4027_/X _4095_/X _5471_/Q vssd1 vssd1 vccd1 vccd1 _4096_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__5788__D _5788_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5150__B _5154_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5244__A3 _2831_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3047_ _3047_/A vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4047__A _5572_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3886__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2790__A _2790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4998_ _4998_/A vssd1 vssd1 vccd1 vccd1 _5631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3949_ _3949_/A _5284_/A vssd1 vssd1 vccd1 vccd1 _3949_/Y sky130_fd_sc_hd__nor2_8
XFILLER_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2766__A1 _5363_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__B1 _3960_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5619_ _5692_/CLK _5619_/D vssd1 vssd1 vccd1 vccd1 _5619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4510__A _4514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3191__A1 input50/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5509__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5659__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input130_A ksc_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5698__D _5698_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2693__B1_N _2692_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4443__A1 _2700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2757__A1 _2592_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2850__D _2850_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5219__C _5219_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output182_A _4010_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3182__A1 _5408_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3681__D _3681_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3036__A _3038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2875__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4793__C _4796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5401__D _5401_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4434__A1 _5376_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4921_ _4921_/A vssd1 vssd1 vccd1 vccd1 _5600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4852_ _4836_/X _4837_/X _3910_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5564_/D sky130_fd_sc_hd__a211o_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _3869_/A _3803_/B vssd1 vssd1 vccd1 vccd1 _3803_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__4198__B1 _4197_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4783_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3945__B1 _3826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3734_ _3961_/A vssd1 vssd1 vccd1 vccd1 _3735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3665_ _3665_/A _4128_/A vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3645__S _3645_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5404_ _5446_/CLK _5404_/D vssd1 vssd1 vccd1 vccd1 _5404_/Q sky130_fd_sc_hd__dfxtp_1
X_2616_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4330__A _4330_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3596_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3613_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5145__B _5154_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2905__D1 _2701_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3173__A1 input47/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5335_ _5741_/CLK _5335_/D vssd1 vssd1 vccd1 vccd1 _5335_/Q sky130_fd_sc_hd__dfxtp_1
X_2547_ _2607_/A vssd1 vssd1 vccd1 vccd1 _2707_/A sky130_fd_sc_hd__buf_2
Xclkbuf_opt_1_1_CLK clkbuf_opt_1_1_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_7_CLK/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5266_ _5266_/A _5266_/B _5266_/C vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__and3_1
XANTENNA__4984__B _4990_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5801__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _3769_/X _3770_/X _4217_/C _4243_/D vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4122__B1 _4109_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2785__A _2785_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5197_ _5197_/A vssd1 vssd1 vccd1 vccd1 _5729_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3476__A2 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5161__A _5161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _5578_/Q vssd1 vssd1 vccd1 vccd1 _4148_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4145_/A _4079_/B _4079_/C vssd1 vssd1 vccd1 vccd1 _4079_/X sky130_fd_sc_hd__and3_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2987__A1 input31/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4505__A _4567_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2739__A1 _2621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5039__C _5039_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5331__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4240__A _4240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__C _4283_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3164__A1 _5405_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4131__B_N _4000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5481__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4113__B1 _4112_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input39_A cpu_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3303__B _5543_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__A1 _2973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__A _4415_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output397_A _3063_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3927__B1 _3925_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3973__B _4079_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3450_ _3281_/A _2899_/A _4674_/C vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2589__B _2589_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3155__A1 input43/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3381_ _3381_/A vssd1 vssd1 vccd1 vccd1 _3381_/X sky130_fd_sc_hd__clkbuf_1
X_5120_ _5120_/A _5130_/B _5236_/A vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__and3_1
XFILLER_83_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4104__B1 _4103_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5051_ _5051_/A vssd1 vssd1 vccd1 vccd1 _5655_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5301__C1 _5278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3458__A2 _2927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4655__A1 _5476_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4002_ _3922_/X _3958_/X _3998_/X _4001_/X vssd1 vssd1 vccd1 vccd1 _4002_/X sky130_fd_sc_hd__o211a_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2666__B1 _4423_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3863__C1 _3862_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5080__A1 _5075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2969__A1 input27/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4904_ _4904_/A vssd1 vssd1 vccd1 vccd1 _5593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3091__A0 _4318_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4325__A _4325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4044__B _4079_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4835_ _4835_/A vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__buf_4
XANTENNA__5354__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _5525_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4591__B1 _4584_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3717_ _2728_/A _3716_/X _5453_/Q vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__a21boi_2
X_4697_ _4697_/A _4707_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__and3_1
XANTENNA__3375__S _3396_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5156__A _5156_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3648_ _4292_/B _5591_/Q _3652_/S vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3146__A1 _5402_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4995__A _5128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3579_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4894__A1 _5590_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5318_ _5741_/CLK _5318_/D vssd1 vssd1 vccd1 vccd1 _5318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4894__B2 _4873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5249_ _2696_/B _2696_/C _4891_/X _5238_/X vssd1 vssd1 vccd1 vccd1 _5755_/D sky130_fd_sc_hd__a211o_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4646__A1 _5468_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2657__B1 _5759_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__B _3134_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5071__A1 _5069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3909__B1 _3831_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4031__C1 _4030_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5066__A _5066_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_22_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4885__A1 _4875_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4637__A1 _5462_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3314__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output312_A _3481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5377__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5062__A1 _4889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2950_ _3157_/A vssd1 vssd1 vccd1 vccd1 _3235_/S sky130_fd_sc_hd__buf_4
XANTENNA__4145__A _4145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4270__C1 _4269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4177__B_N _4083_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2820__B1 _2819_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2881_ _4295_/B vssd1 vssd1 vccd1 vccd1 _2882_/A sky130_fd_sc_hd__buf_4
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4620_ _4645_/A vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _5422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3502_ _3504_/A _5646_/Q vssd1 vssd1 vccd1 vccd1 _3503_/A sky130_fd_sc_hd__and2_1
X_4482_ _4482_/A vssd1 vssd1 vccd1 vccd1 _5395_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5117__A2 _2899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3128__A1 _5399_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3433_ _3445_/A _3433_/B _4749_/C vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__and3_1
XFILLER_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3679__A2 _4746_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4030__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3364_ _4322_/B _5499_/Q _3364_/S vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__mux2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5099_/X _5094_/X _5087_/X _5102_/X _4159_/B vssd1 vssd1 vccd1 vccd1 _5683_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3295_ _3303_/A _5539_/Q vssd1 vssd1 vccd1 vccd1 _3296_/A sky130_fd_sc_hd__and2_1
XFILLER_100_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__clkbuf_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3878__B _4283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2782__B _2782_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5796__D _5796_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4055__A _4055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4261__C1 _4153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2811__B1 _2690_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4205__D _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4818_ _4818_/A vssd1 vssd1 vccd1 vccd1 _5549_/D sky130_fd_sc_hd__clkbuf_1
X_5798_ _5798_/CLK _5798_/D vssd1 vssd1 vccd1 vccd1 _5798_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4749_/A _4763_/B _4749_/C vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__or3_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5108__A2 _4837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5036__D _5043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4867__A1 _4859_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput103 gpio_dat_i[7] vssd1 vssd1 vccd1 vccd1 _3907_/C sky130_fd_sc_hd__clkbuf_1
Xinput114 ksc_dat_i[14] vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput125 ksc_dat_i[24] vssd1 vssd1 vccd1 vccd1 _4184_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 ksc_dat_i[5] vssd1 vssd1 vccd1 vccd1 _5073_/B2 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4619__A1 _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput147 spi_dat_i[12] vssd1 vssd1 vccd1 vccd1 _3996_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4108__A2_N _5680_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput158 spi_dat_i[22] vssd1 vssd1 vccd1 vccd1 _4161_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput169 spi_dat_i[3] vssd1 vssd1 vccd1 vccd1 _3820_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5292__A1 _5783_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5292__B2 _4034_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2973__A _3042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3842__A2 _3804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2802__B1 _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3699__A_N _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3309__A _3309_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4131__C _4131_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output262_A _3430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4858__A1 _3960_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4858__B2 _4857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3970__C _4143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2869__B1 _5058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2867__B _3697_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3044__A _3849_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ _4312_/B _5391_/Q _3248_/S vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4086__A2 _3906_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5283__A1 _5777_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5283__B2 _3928_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3979__A _3979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5035__A1 _5646_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5035__B2 _5034_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3982_ _3977_/X _3978_/X _3979_/X _3981_/X _3908_/X vssd1 vssd1 vccd1 vccd1 _3982_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3210__C _4526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3597__A1 _5612_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2933_ _4423_/C _4423_/B _2689_/Y _2932_/Y vssd1 vssd1 vccd1 vccd1 _2937_/B sky130_fd_sc_hd__a211oi_2
X_5721_ _5741_/CLK _5721_/D vssd1 vssd1 vccd1 vccd1 _5721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5652_ _5659_/CLK _5652_/D vssd1 vssd1 vccd1 vccd1 _5652_/Q sky130_fd_sc_hd__dfxtp_1
X_2864_ _2864_/A _2864_/B _4405_/A vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__nand3_2
X_4603_ _5444_/Q _4589_/X _4584_/X _4590_/X _4598_/X vssd1 vssd1 vccd1 vccd1 _5444_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4322__B _4322_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5583_ _5694_/CLK _5583_/D vssd1 vssd1 vccd1 vccd1 _5583_/Q sky130_fd_sc_hd__dfxtp_1
X_2795_ _2795_/A _2864_/A _2864_/B _2795_/D vssd1 vssd1 vccd1 vccd1 _2796_/C sky130_fd_sc_hd__nand4_1
X_4534_ _4538_/A _4550_/B _4534_/C vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__or3_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4041__C _4143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _5389_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4976__C _4976_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4849__A1 _3662_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3416_ _3429_/A _3416_/B _4737_/A vssd1 vssd1 vccd1 vccd1 _3417_/A sky130_fd_sc_hd__and3_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4396_ _4396_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__and2_1
XFILLER_63_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5542__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3347_ _4310_/A _5494_/Q _3441_/S vssd1 vssd1 vccd1 vccd1 _4688_/C sky130_fd_sc_hd__mux2_1
XFILLER_24_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5259__D1 _4429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3316_/A vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__buf_2
XANTENNA__4992__B _4997_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5021_/A _5639_/Q _5017_/C _5021_/D vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__and4_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3401__B _3416_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4234__C1 _4233_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4785__B1 _3723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4513__A _4513_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3129__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5047__C _5056_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2968__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input160_A spi_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2687__B _2831_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input21_A cpu_adr_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__A2 _3915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3276__B1 _4778_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4423__A _4431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5415__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3684__D _5094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3039__A _3039_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2580_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2848_/B sky130_fd_sc_hd__clkbuf_4
Xoutput407 _3227_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput418 _3241_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__3751__A1 _5662_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2878__A _2878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5565__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__B2 _5065_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3473__S _3652_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4796__C _4796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4250_ _4250_/A vssd1 vssd1 vccd1 vccd1 _4250_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3201_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3201_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4181_ _4042_/X _4175_/Y _4180_/Y _4153_/X vssd1 vssd1 vccd1 vccd1 _4181_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5404__D _5404_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3132_ _5162_/C _5330_/Q _3132_/S vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__mux2_8
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3205__C _4524_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _3063_/A vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3502__A _3504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3221__B _3221_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3965_ _5779_/Q _3915_/X _3953_/X _3964_/Y vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__o22ai_4
XANTENNA__3648__S _3652_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5704_ _5766_/CLK _5704_/D vssd1 vssd1 vccd1 vccd1 _5704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2916_ _2916_/A _2916_/B _2916_/C _2929_/C vssd1 vssd1 vccd1 vccd1 _2917_/C sky130_fd_sc_hd__nand4_1
XANTENNA__4333__A _4333_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3896_ _5775_/Q _3690_/X _3886_/X _3895_/Y vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__o22ai_4
XANTENNA__2793__A2 _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5148__B _5167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5635_ _5635_/CLK _5635_/D vssd1 vssd1 vccd1 vccd1 _5635_/Q sky130_fd_sc_hd__dfxtp_1
X_2847_ _2809_/X _2750_/X _5360_/Q vssd1 vssd1 vccd1 vccd1 _2850_/C sky130_fd_sc_hd__o21ai_1
XFILLER_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5566_ _5586_/CLK _5566_/D vssd1 vssd1 vccd1 vccd1 _5566_/Q sky130_fd_sc_hd__dfxtp_1
X_2778_ _4098_/A vssd1 vssd1 vccd1 vccd1 _2778_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4517_ _4517_/A _4526_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__and3_1
XANTENNA__2788__A _2788_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5497_ _5538_/CLK _5497_/D vssd1 vssd1 vccd1 vccd1 _5497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3383__S _3396_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5164__A _5212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4448_ _5204_/A vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__buf_2
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4431_/A vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__buf_2
XANTENNA__5314__D _5314_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2702__C1 _2932_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3732__B_N _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5247__A1 _2715_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4508__A _4508_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3412__A _3412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5438__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4222__A2 _4091_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5058__B _5058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2784__A2 _2671_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5588__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3733__A1 _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input69_A cpu_sel_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2698__A _2698_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3306__B _5544_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2848__D _2848_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3249__B1 _4454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4418__A _4418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output225_A _3311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3322__A _3322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2864__C _4405_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3917__A1_N _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4137__B _4137_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2880__B _2925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4153__A _4153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3750_ _3846_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__buf_2
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _5764_/Q _2683_/X _2698_/Y _2699_/X _2700_/X vssd1 vssd1 vccd1 vccd1 _2701_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _3742_/A _3681_/B _3681_/C _3681_/D vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__nand4_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5420_ _5435_/CLK _5420_/D vssd1 vssd1 vccd1 vccd1 _5420_/Q sky130_fd_sc_hd__dfxtp_1
X_2632_ _5372_/Q vssd1 vssd1 vccd1 vccd1 _2632_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput204 _3843_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[3] sky130_fd_sc_hd__buf_2
X_5351_ _5737_/CLK _5351_/D vssd1 vssd1 vccd1 vccd1 _5351_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput215 _3291_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[13] sky130_fd_sc_hd__buf_2
X_2563_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2622_/A sky130_fd_sc_hd__buf_2
Xoutput226 _3313_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[23] sky130_fd_sc_hd__buf_2
XFILLER_86_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput237 _3270_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput248 _3385_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[13] sky130_fd_sc_hd__buf_2
X_4302_ _4302_/A vssd1 vssd1 vccd1 vccd1 _5316_/D sky130_fd_sc_hd__clkbuf_1
Xoutput259 _3421_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[23] sky130_fd_sc_hd__buf_2
X_5282_ _5282_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5776_/D sky130_fd_sc_hd__nand2_1
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3216__B _3221_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4233_ _4230_/Y _4115_/X _4232_/Y vssd1 vssd1 vccd1 vccd1 _4233_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4164_ _3735_/A _4003_/A _5579_/Q vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__o21a_2
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5229__A1 _2836_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3115_ _5154_/A _5327_/Q _3162_/S vssd1 vssd1 vccd1 vccd1 _4327_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4328__A _4328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4095_ _4110_/A vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3232__A _3232_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3062_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5150__C _5160_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3886__B _3886_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4997_ _4997_/A _4997_/B _4997_/C vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__and3_1
XFILLER_36_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5159__A _5183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5730__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3948_ _5778_/Q _3804_/X _3936_/X _3947_/Y vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__o22ai_4
XFILLER_36_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2766__A2 _2696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__A1 _3720_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__B2 _3962_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4998__A _4998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3879_ _5458_/Q _4444_/A _3878_/X vssd1 vssd1 vccd1 vccd1 _3879_/Y sky130_fd_sc_hd__a21oi_4
X_5618_ _5692_/CLK _5618_/D vssd1 vssd1 vccd1 vccd1 _5618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3701__A2_N _5661_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5549_ _5555_/CLK _5549_/D vssd1 vssd1 vccd1 vccd1 _5549_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4510__B _4524_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3407__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4238__A _4238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__A _3142_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input123_A ksc_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4443__A2 _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3651__B1 _4901_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__A _5096_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2757__A2 _2790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4701__A _4701_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3317__A _3325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3036__B _5448_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output342_A _3556_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5603__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4148__A _5578_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2693__A1 _2675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3052__A _3163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4434__A2 _4429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3987__A _4036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5092__C1 _4058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5753__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2891__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4920_ _4938_/A _4938_/B _4920_/C vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__or3_1
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3642__A0 _4371_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4851_ _3892_/X _3893_/X _4832_/X _4833_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _5563_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3198__S _3219_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3802_ _5771_/Q _3690_/X _3792_/X _3801_/Y vssd1 vssd1 vccd1 vccd1 _3803_/B sky130_fd_sc_hd__o22ai_4
XANTENNA__4198__B2 _4141_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4782_ _4804_/A vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3902__A_N _3817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3945__A1 _3940_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3733_ _3277_/A _3723_/X _3725_/X _3732_/X vssd1 vssd1 vccd1 vccd1 _3733_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4611__A _4611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3664_ _3664_/A vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__buf_2
X_5403_ _5446_/CLK _5403_/D vssd1 vssd1 vccd1 vccd1 _5403_/Q sky130_fd_sc_hd__dfxtp_1
X_2615_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__buf_4
X_3595_ _3595_/A vssd1 vssd1 vccd1 vccd1 _3595_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3227__A _3227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2905__C1 _2932_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3809__A1_N _3806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5145__C _5160_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2546_ _5767_/Q vssd1 vssd1 vccd1 vccd1 _2607_/A sky130_fd_sc_hd__buf_4
X_5334_ _5741_/CLK _5334_/D vssd1 vssd1 vccd1 vccd1 _5334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5265_ _5265_/A vssd1 vssd1 vccd1 vccd1 _5766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4984__C _4984_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4122__A1 _5788_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__B2 _4121_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4216_ _4216_/A1 _4449_/A _3994_/A _4215_/Y vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__a31oi_4
X_5196_ _5200_/A _5215_/B _5196_/C vssd1 vssd1 vccd1 vccd1 _5197_/A sky130_fd_sc_hd__or3_1
XFILLER_96_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5799__D _5799_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4147_/A vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4058__A _4127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3881__B1 _3877_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4421__C_N _2932_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4075_/X _4076_/X _4078_/C _4201_/D vssd1 vssd1 vccd1 vccd1 _4079_/C sky130_fd_sc_hd__and4bb_1
XFILLER_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3897__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5083__C1 _3970_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3029_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3038_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3633__A0 _4364_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_2_0_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2739__A2 _2696_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5039__D _5043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__A _4521_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4240__B _4240_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__D _3782_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3137__A _3250_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5626__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4113__A1 _5472_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2695__B _2695_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5776__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5502__D _5502_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5074__C1 _3886_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2978__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__B _4415_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3927__A1 _3720_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output292_A _3505_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3927__B2 _3926_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4431__A _4431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3973__C _3973_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3047__A _3047_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2589__C _2589_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4888__C1 _4848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3380_ _3393_/A _3380_/B _4712_/A vssd1 vssd1 vccd1 vccd1 _3381_/A sky130_fd_sc_hd__and3_1
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5050_ _5056_/A _5655_/Q _5056_/C _5056_/D vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__and4_1
XFILLER_65_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4104__A1 _4059_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5301__B1 _4159_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4001_ _3999_/X _4000_/X _4001_/C _4063_/D vssd1 vssd1 vccd1 vccd1 _4001_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4655__A2 _4652_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2666__A1 _5371_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5412__D _5412_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3863__B1 _3768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5065__C1 _5111_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3510__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5080__A2 _4890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4903_ _4903_/A _4915_/B _4915_/C vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__and3_1
XANTENNA__3091__A1 _5393_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4834_ _3733_/X _3738_/X _4832_/X _4833_/X _4630_/X vssd1 vssd1 vccd1 vccd1 _5557_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4044__C _4044_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4765_ _4765_/A _4778_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__and3_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4591__A1 _5438_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4341__A _4341_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3716_ _4110_/A vssd1 vssd1 vccd1 vccd1 _3716_/X sky130_fd_sc_hd__buf_2
XANTENNA__5649__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4591__B2 _4590_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4696_ _4778_/C vssd1 vssd1 vccd1 vccd1 _4716_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4879__C1 _4865_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3578_ _3578_/A vssd1 vssd1 vccd1 vccd1 _3578_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4995__B _5005_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4894__A2 _4688_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _5766_/CLK _5317_/D vssd1 vssd1 vccd1 vccd1 _5317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2796__A _2796_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5799__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5172__A _5176_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5248_ _5754_/Q _5234_/X _2831_/Y _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5754_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4646__A2 _4639_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2657__A1 _2695_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5322__D _5322_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5179_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5722_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3854__B1 _3669_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__C _4487_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4516__A _4595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3420__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5071__A2 _4890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3909__A1 _3829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__B1 _3998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input51_A cpu_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4885__A2 _4876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4637__A2 _4623_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3314__B _5548_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output305_A _3529_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4426__A _4426_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3330__A _3330_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5062__A2 _5060_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4270__B1 _3831_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4145__B _4228_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2820__A1 _5762_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2880_ _2909_/A _2925_/A _2887_/C _2925_/B vssd1 vssd1 vccd1 vccd1 _4295_/B sky130_fd_sc_hd__and4_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4550_ _4674_/A _4550_/B _4550_/C vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__or3_1
XANTENNA__4253__A_N _4075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3501_ _3501_/A vssd1 vssd1 vccd1 vccd1 _3501_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5407__D _5407_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4481_ _4481_/A _4500_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__and3_1
X_3432_ _4364_/A _5518_/Q _3432_/S vssd1 vssd1 vccd1 vccd1 _4749_/C sky130_fd_sc_hd__mux2_1
XFILLER_83_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3363_ _3418_/A vssd1 vssd1 vccd1 vccd1 _3380_/B sky130_fd_sc_hd__clkbuf_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3505__A _3505_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5102_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5102_/X sky130_fd_sc_hd__buf_2
X_3294_ _3316_/A vssd1 vssd1 vccd1 vccd1 _3303_/A sky130_fd_sc_hd__clkbuf_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4089__B1 _4073_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__C1 _5285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__clkbuf_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5038__C1 _5023_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5321__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4336__A _4336_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__C _4283_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2782__C _2782_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4261__B1 _4260_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2811__A1 _2809_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5471__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4817_ _4821_/A _5549_/Q _4817_/C vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__and3_1
XANTENNA__3386__S _3400_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5797_ _5802_/CLK _5797_/D vssd1 vssd1 vccd1 vccd1 _5797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5167__A _5176_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4071__A _4071_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4748_ _4748_/A vssd1 vssd1 vccd1 vccd1 _5517_/D sky130_fd_sc_hd__clkbuf_1
X_4679_ _4699_/A _4688_/B _4679_/C vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__or3_1
XANTENNA__5317__D _5317_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5108__A3 _4872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4867__A2 _4860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput104 gpio_dat_i[8] vssd1 vssd1 vccd1 vccd1 _3924_/C sky130_fd_sc_hd__buf_2
XFILLER_66_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput115 ksc_dat_i[15] vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput126 ksc_dat_i[25] vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4619__A2 _3857_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput137 ksc_dat_i[6] vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3134__B _3134_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput148 spi_dat_i[13] vssd1 vssd1 vccd1 vccd1 _4018_/D sky130_fd_sc_hd__clkbuf_2
Xinput159 spi_dat_i[23] vssd1 vssd1 vccd1 vccd1 _4173_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5292__A2 _5289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2802__A1 _2778_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input99_A gpio_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4004__B1 _5569_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5805__A _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4131__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4858__A2 _3962_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3970__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output255_A _3340_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2869__A1 _2859_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3325__A _3325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output422_A _5807_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5283__A2 _5269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4144__B_N _4076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4156__A _4195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3060__A _3163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5035__A2 _5033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5494__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3832_/X _3833_/X _3981_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _3981_/X sky130_fd_sc_hd__and4bb_1
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5720_ _5741_/CLK _5720_/D vssd1 vssd1 vccd1 vccd1 _5720_/Q sky130_fd_sc_hd__dfxtp_1
X_2932_ _2932_/A _2932_/B _2932_/C _2932_/D vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__nand4_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5651_ _5659_/CLK _5651_/D vssd1 vssd1 vccd1 vccd1 _5651_/Q sky130_fd_sc_hd__dfxtp_1
X_2863_ _2916_/A _2916_/B _2916_/C _2929_/C vssd1 vssd1 vccd1 vccd1 _2866_/C sky130_fd_sc_hd__and4_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4602_ _4602_/A vssd1 vssd1 vccd1 vccd1 _5443_/D sky130_fd_sc_hd__clkbuf_1
X_5582_ _5586_/CLK _5582_/D vssd1 vssd1 vccd1 vccd1 _5582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2794_ _2794_/A _2852_/C _2794_/C vssd1 vssd1 vccd1 vccd1 _2796_/B sky130_fd_sc_hd__nand3_1
X_4533_ _4533_/A vssd1 vssd1 vccd1 vccd1 _5415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4041__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _4464_/A _4475_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__and3_1
XANTENNA__4849__A2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3415_ _4353_/B _5513_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _5356_/D sky130_fd_sc_hd__clkbuf_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3346_ _3445_/B vssd1 vssd1 vccd1 vccd1 _3361_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__C1 _4848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4149__A_N _4082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3277_/A vssd1 vssd1 vccd1 vccd1 _3316_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__B1 _3807_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4992__C _4997_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5638_/Q _5010_/X _5806_/A _5011_/X _4823_/X vssd1 vssd1 vccd1 vccd1 _5638_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5600__D _5600_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_21_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3401__C _4726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__B1 _3758_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4785__A1 _3316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3129__B _3134_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5047__D _5056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5367__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2687__C _2813_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input153_A spi_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2720__B1 _5754_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3276__A1 _3267_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A cpu_adr_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5510__D _5510_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4225__B1 _4224_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4704__A _4917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3984__C1 _3983_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4423__B _4423_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output372_A _3035_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput408 _3069_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__3981__C _3981_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput419 _3245_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__3751__A2 _5002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2878__B _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3055__A _3055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3200_ _3210_/A _3221_/B _4522_/A vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__and3_1
XFILLER_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4180_ _4147_/X _4046_/X _3758_/A _4179_/Y vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__2894__A _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3131_ _5715_/Q input39/X _3168_/S vssd1 vssd1 vccd1 vccd1 _5162_/C sky130_fd_sc_hd__mux2_1
XFILLER_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5270__A _5270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3062_ _3062_/A _3073_/B _4460_/C vssd1 vssd1 vccd1 vccd1 _3063_/A sky130_fd_sc_hd__and3_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3502__B _5646_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5420__D _5420_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3221__C _4532_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4216__B1 _4215_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4614__A _4652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3964_ _3887_/X _4638_/B _3963_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _3964_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5703_ _5765_/CLK _5703_/D vssd1 vssd1 vccd1 vccd1 _5703_/Q sky130_fd_sc_hd__dfxtp_1
X_2915_ _2895_/X _2899_/X _4761_/A vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4333__B _4333_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3895_ _3887_/X _4634_/B _3894_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _3895_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5634_ _5694_/CLK _5634_/D vssd1 vssd1 vccd1 vccd1 _5634_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5148__C _5148_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2846_ _2806_/X _2699_/X _5363_/Q vssd1 vssd1 vccd1 vccd1 _2846_/Y sky130_fd_sc_hd__a21oi_1
X_5565_ _5802_/CLK _5565_/D vssd1 vssd1 vccd1 vccd1 _5565_/Q sky130_fd_sc_hd__dfxtp_1
X_2777_ _5556_/Q vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__clkbuf_2
X_4516_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4536_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3891__C _3891_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5496_ _5538_/CLK _5496_/D vssd1 vssd1 vccd1 vccd1 _5496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2788__B _2788_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4447_ _4466_/A vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__buf_12
XFILLER_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__C1 _4151_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4378_ _4378_/A vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2702__B1 _2932_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A cpu_adr_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3329_ _3329_/A _5555_/Q vssd1 vssd1 vccd1 vccd1 _3330_/A sky130_fd_sc_hd__and2_1
XFILLER_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5180__A _5204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__A2 _5227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4508__B _4526_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3412__B _3416_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5330__D _5330_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4227__C _4227_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4207__B1 _4206_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__A _4538_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2769__B1 _5556_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2784__A3 _2574_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5058__C _5235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3733__A2 _3723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2698__B _2831_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5505__D _5505_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5090__A _5090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3603__A _3622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3249__A1 _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output218_A _3298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2880__C _2887_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5532__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2700_ _2806_/A vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__clkbuf_4
X_3680_ _3680_/A _3757_/A _3682_/A vssd1 vssd1 vccd1 vccd1 _3681_/D sky130_fd_sc_hd__nand3_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _2878_/A _2909_/A _2929_/A vssd1 vssd1 vccd1 vccd1 _2631_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__5265__A _5265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5350_ _5737_/CLK _5350_/D vssd1 vssd1 vccd1 vccd1 _5350_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput205 _3869_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[4] sky130_fd_sc_hd__buf_2
X_2562_ _2675_/A _2559_/X _2560_/Y _2561_/Y vssd1 vssd1 vccd1 vccd1 _2589_/B sky130_fd_sc_hd__o211a_1
Xoutput216 _3293_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[14] sky130_fd_sc_hd__buf_2
XANTENNA__5682__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput227 _3315_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__4093__A2_N _5679_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput238 _3272_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[5] sky130_fd_sc_hd__buf_2
X_4301_ _4301_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__or2_1
Xoutput249 _3388_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5281_ _5775_/Q _5269_/X _3886_/X _3895_/Y _5310_/B vssd1 vssd1 vccd1 vccd1 _5775_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5415__D _5415_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4134__C1 _4005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3216__C _4529_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4232_ _3763_/A _3766_/A _3768_/A _4231_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4232_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4609__A _4609_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4163_ _4098_/X _3958_/A _4781_/A _4162_/X vssd1 vssd1 vccd1 vccd1 _4163_/X sky130_fd_sc_hd__o211a_1
XFILLER_99_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3513__A _3515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5229__A2 _5227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3114_ _3174_/A vssd1 vssd1 vccd1 vccd1 _3162_/S sky130_fd_sc_hd__buf_4
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4094_ _4127_/A _4094_/B _4159_/C _4214_/D vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__and4_2
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3045_ _3878_/A vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__buf_2
XANTENNA__3981__A_N _3832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3886__C _3993_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4344__A _4344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _5630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3947_ _3813_/X _3939_/Y _3945_/Y _3946_/X vssd1 vssd1 vccd1 vccd1 _3947_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3963__A2 _3890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3878_ _3878_/A _4283_/B _4283_/C _3878_/D vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__and4_2
X_5617_ _5692_/CLK _5617_/D vssd1 vssd1 vccd1 vccd1 _5617_/Q sky130_fd_sc_hd__dfxtp_1
X_2829_ _5369_/Q vssd1 vssd1 vccd1 vccd1 _2829_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2799__A _5590_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3176__A0 _4349_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5175__A _5175_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5548_ _5555_/CLK _5548_/D vssd1 vssd1 vccd1 vccd1 _5548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4510__C _4510_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5325__D _5325_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5479_ _5482_/CLK _5479_/D vssd1 vssd1 vccd1 vccd1 _5479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4519__A _4678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3423__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5405__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4205__B_N _4083_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A ksc_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A1 _3482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5555__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__S _3597_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A _4254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input81_A gpio_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4701__B _4707_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3317__B _5549_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output335_A _3638_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4429__A _5264_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__A _3453_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2693__A2 _2750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4419__B1 _4402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5092__B1 _5084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3987__B _5288_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A1 _5625_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4836_/X _4837_/X _3875_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5562_/D sky130_fd_sc_hd__a211o_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _3707_/X _4626_/B _3800_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _3801_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4804_/A sky130_fd_sc_hd__buf_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3732_ _3727_/X _3729_/X _3732_/C _3978_/A vssd1 vssd1 vccd1 vccd1 _3732_/X sky130_fd_sc_hd__and4bb_1
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3945__A2 _3825_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4611__B _5449_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3663_ _3823_/A _3755_/A _3678_/A _3662_/Y _3683_/A vssd1 vssd1 vccd1 vccd1 _3742_/A
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3158__A0 _4342_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3508__A _3508_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5402_ _5731_/CLK _5402_/D vssd1 vssd1 vccd1 vccd1 _5402_/Q sky130_fd_sc_hd__dfxtp_1
X_2614_ _2614_/A vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__inv_2
X_3594_ _3594_/A _3601_/B _4949_/A vssd1 vssd1 vccd1 vccd1 _3595_/A sky130_fd_sc_hd__and3_1
XANTENNA__2905__B1 _2932_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5333_ _5695_/CLK _5333_/D vssd1 vssd1 vccd1 vccd1 _5333_/Q sky130_fd_sc_hd__dfxtp_1
X_2545_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5428__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5264_ _5264_/A _5266_/B _5264_/C vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__and3_1
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4215_ _3878_/A _4095_/X _5479_/Q vssd1 vssd1 vccd1 vccd1 _4215_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_29_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4122__A2 _4070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4339__A _4339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2669__C1 _2637_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5195_ _5195_/A vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _5474_/Q _4074_/X _4145_/X vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4058__B _4058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3881__A1 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5578__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3881__B2 _3880_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4253_/D vssd1 vssd1 vccd1 vccd1 _4201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5083__B1 _5076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3897__B _3897_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3028_ _3028_/A vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3633__A1 _5622_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3389__S _3396_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4074__A _4074_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _4979_/A vssd1 vssd1 vccd1 vccd1 _5623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4594__C1 _4576_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4802__A _4802_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2739__A3 _2696_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3149__A0 _5718_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3418__A _3418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4240__C _4240_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4113__A2 _4074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4249__A _4263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3153__A _3153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2695__C _2695_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2992__A _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5074__B1 _5061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__C1 _2606_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__C _4439_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4585__C1 _4576_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4712__A _4712_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3927__A2 _3890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4431__B _4431_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output285_A _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3328__A _3328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4888__B1 _4271_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2589__D _4411_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5301__A1 _5791_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4104__A2 _4649_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5301__B2 _4166_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4159__A _4240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5720__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3063__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _4000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3863__A1 _3763_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2666__A2 _2611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3998__A _3998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5065__B1 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4273__D1 _3866_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _4902_/A vssd1 vssd1 vccd1 vccd1 _5592_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5080__A3 _5070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ _5087_/A vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__A0 _4331_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4622__A _4638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4764_ _4764_/A vssd1 vssd1 vccd1 vccd1 _5524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _3850_/A vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4591__A2 _4589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4695_ _4695_/A vssd1 vssd1 vccd1 vccd1 _5496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3646_ _3646_/A _4988_/B _4984_/C vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__and3_1
XANTENNA__4879__B1 _4872_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3577_ _3577_/A _3584_/B _4934_/C vssd1 vssd1 vccd1 vccd1 _3578_/A sky130_fd_sc_hd__and3_1
XANTENNA__3551__A0 _4312_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4995__C _4995_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5316_ _5741_/CLK _5316_/D vssd1 vssd1 vccd1 vccd1 _5316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2796__B _2796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5172__B _5191_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5247_ _2715_/Y _5227_/X _2716_/Y _4848_/A _4429_/X vssd1 vssd1 vccd1 vccd1 _5753_/D
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__4069__A _4123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5603__D _5603_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5178_ _5178_/A _5178_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__and3_1
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2657__A2 _2695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3854__A1 _2845_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4129_ _4027_/X _4095_/X _5473_/Q vssd1 vssd1 vccd1 vccd1 _4129_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3420__B _3433_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5071__A3 _5070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2814__C1 _2606_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4532__A _4532_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3909__A2 _3830_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__A1 _3922_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3148__A _3148_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5743__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input44_A cpu_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5513__D _5513_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4707__A _4707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3611__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output200_A _4263_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5062__A3 _4847_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__A1 _3829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4145__C _4145_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2820__A2 _2577_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4442__A _4442_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3058__A _3144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3500_ _3504_/A _5645_/Q vssd1 vssd1 vccd1 vccd1 _3501_/A sky130_fd_sc_hd__and2_1
XFILLER_89_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4480_ _5228_/A vssd1 vssd1 vccd1 vccd1 _4500_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3431_ _3431_/A vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2897__A _2925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5273__A _5299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3362_ _3362_/A vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__clkbuf_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5096_/X _5089_/X _5090_/X _5097_/X _4143_/B vssd1 vssd1 vccd1 vccd1 _5682_/D
+ sky130_fd_sc_hd__a311o_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3293_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3293_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5423__D _5423_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4089__A1 _5786_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__B1 _3953_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4089__B2 _4088_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5645_/D sky130_fd_sc_hd__clkbuf_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4617__A _4617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3521__A _3521_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5038__B1 _5029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3878__D _3878_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2782__D _2782_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4261__A1 _3792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5616__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2811__A2 _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4816_ _5548_/Q _4803_/X _4798_/X _4804_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5548_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4352__A _4352_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4078__A_N _4075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5796_ _5798_/CLK _5796_/D vssd1 vssd1 vccd1 vccd1 _5796_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5167__B _5167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4747_ _4747_/A _4756_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__and3_1
XANTENNA__5766__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4678_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3629_ _4362_/B _5621_/Q _3636_/S vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5183__A _5183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2600__A _2622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput105 gpio_dat_i[9] vssd1 vssd1 vccd1 vccd1 _3942_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5333__D _5333_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput116 ksc_dat_i[16] vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput127 ksc_dat_i[26] vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput138 ksc_dat_i[7] vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3134__C _4494_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput149 spi_dat_i[14] vssd1 vssd1 vccd1 vccd1 _4029_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4527__A _4527_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3431__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2802__A2 _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4004__A1 _3961_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5508__D _5508_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3606__A _3613_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2869__A2 _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3325__B _5553_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2723__D1 _2787_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output248_A _3385_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4437__A _4441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output415_A _3100_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3341__A _4830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5639__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4156__B _5300_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _4149_/D sky130_fd_sc_hd__clkbuf_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2931_ _5266_/C _2676_/X _5372_/Q vssd1 vssd1 vccd1 vccd1 _2932_/A sky130_fd_sc_hd__o21ai_1
XFILLER_91_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5789__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5268__A _5268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5650_ _5659_/CLK _5650_/D vssd1 vssd1 vccd1 vccd1 _5650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4172__A _4252_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2862_ _2809_/A _2559_/X _2861_/Y _2859_/Y vssd1 vssd1 vccd1 vccd1 _2929_/C sky130_fd_sc_hd__o211a_1
X_4601_ _4611_/A _5443_/Q _4604_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__and4_1
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5581_ _5589_/CLK _5581_/D vssd1 vssd1 vccd1 vccd1 _5581_/Q sky130_fd_sc_hd__dfxtp_1
X_2793_ _5362_/Q _2903_/A _2792_/Y vssd1 vssd1 vccd1 vccd1 _2852_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__5418__D _5418_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4532_ _4532_/A _4556_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__and3_1
XANTENNA__4900__A _4968_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4463_ _4652_/A vssd1 vssd1 vccd1 vccd1 _4485_/C sky130_fd_sc_hd__buf_2
XANTENNA__3516__A _3516_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3414_ _3431_/A vssd1 vssd1 vccd1 vccd1 _3429_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__4849__A3 _4847_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4394_ _4394_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__or2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3345_/A vssd1 vssd1 vccd1 vccd1 _3445_/B sky130_fd_sc_hd__buf_2
XFILLER_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__B1 _2641_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3267_/X _3268_/X _4778_/A vssd1 vssd1 vccd1 vccd1 _3276_/X sky130_fd_sc_hd__o21a_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__B2 _3808_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4347__A _4347_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4234__A1 _4147_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4785__A2 _4804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5178__A _5178_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4082__A _4082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5328__D _5328_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5779_ _5802_/CLK _5779_/D vssd1 vssd1 vccd1 vccd1 _5779_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3745__B1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3129__C _4491_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3426__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_22_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5800_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2687__D _2831_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4170__B1 _4169_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2720__A1 _2593_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input146_A spi_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3276__A2 _3268_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4243__A_N _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4225__B2 _4141_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3984__B1 _3975_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4423__C _4423_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output198_A _4237_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4720__A _4720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput409 _3232_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__3981__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output365_A _3020_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3336__A _3336_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4161__B1 _4160_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4111__B_N _4076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3130_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5461__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5270__B _5270_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3061_ _4306_/A _5388_/Q _3230_/S vssd1 vssd1 vccd1 vccd1 _4460_/C sky130_fd_sc_hd__mux2_1
XFILLER_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5110__C1 _4252_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5701__D _5701_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4216__A1 _4216_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _3720_/X _3890_/X _3960_/X _3962_/X _3740_/X vssd1 vssd1 vccd1 vccd1 _3963_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4614__B _5451_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2914_ _3418_/A vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__clkbuf_2
X_5702_ _5766_/CLK _5702_/D vssd1 vssd1 vccd1 vccd1 _5702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3894_ _3720_/X _3890_/X _3892_/X _3893_/X _3740_/X vssd1 vssd1 vccd1 vccd1 _3894_/Y
+ sky130_fd_sc_hd__o221ai_4
X_5633_ _5641_/CLK _5633_/D vssd1 vssd1 vccd1 vccd1 _5633_/Q sky130_fd_sc_hd__dfxtp_1
X_2845_ _5486_/Q vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__buf_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4630__A _4848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5564_ _5586_/CLK _5564_/D vssd1 vssd1 vccd1 vccd1 _5564_/Q sky130_fd_sc_hd__dfxtp_1
X_2776_ _5268_/B vssd1 vssd1 vccd1 vccd1 _2776_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4515_ _4515_/A vssd1 vssd1 vccd1 vccd1 _5408_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3891__D _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4116__A_N _4082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5495_ _5538_/CLK _5495_/D vssd1 vssd1 vccd1 vccd1 _5495_/Q sky130_fd_sc_hd__dfxtp_1
X_4446_ _4446_/A vssd1 vssd1 vccd1 vccd1 _5383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4152__B1 _3975_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4377_ _5264_/C vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2702__A1 _2690_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3328_ _3328_/A vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__clkbuf_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5101__C1 _4143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3259_ _4383_/B _5525_/Q _4803_/A vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5611__D _5611_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__A _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4508__C _4512_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3412__C _4733_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3663__C1 _3683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4227__D _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4805__A _4823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4207__A1 _4204_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4524__B _4524_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2769__A1 _2877_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4243__C _4243_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5334__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3718__B1 _3717_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4540__A _4567_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2698__C _2813_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5484__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2995__A _2995_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3590__S _3597_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3249__A2 _2882_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5521__D _5521_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4715__A _4715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2880__D _2925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4450__A _4558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2630_ _4405_/A _2864_/A _2864_/B vssd1 vssd1 vccd1 vccd1 _2929_/A sky130_fd_sc_hd__and3_1
X_2561_ _5452_/Q vssd1 vssd1 vccd1 vccd1 _2561_/Y sky130_fd_sc_hd__inv_2
Xoutput206 _3882_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput217 _3296_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[15] sky130_fd_sc_hd__buf_2
X_4300_ _4300_/A vssd1 vssd1 vccd1 vccd1 _5315_/D sky130_fd_sc_hd__clkbuf_1
Xoutput228 _3318_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[25] sky130_fd_sc_hd__buf_2
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4289__A_N _4295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput239 _3274_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[6] sky130_fd_sc_hd__buf_2
X_5280_ _5280_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5774_/D sky130_fd_sc_hd__nand2_1
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _3999_/A _4000_/A _4231_/C _4257_/D vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__and4bb_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4134__B1 _4132_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4162_ _3769_/X _3770_/X _4162_/C _4243_/D vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__and4bb_1
XFILLER_64_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3513__B _5651_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3113_ _5712_/Q input36/X _3126_/S vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5431__D _5431_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4093_ _3989_/X _5679_/Q _4092_/Y _3991_/X vssd1 vssd1 vccd1 vccd1 _4094_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3044_ _3849_/A vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3886__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4344__B _4344_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5357__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4995_ _5128_/A _5005_/B _4995_/C vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__or3_1
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3948__B1 _3936_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3946_ _4153_/A vssd1 vssd1 vccd1 vccd1 _3946_/X sky130_fd_sc_hd__buf_2
XANTENNA__4063__C _4063_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2620__B1 _2619_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3877_ _3871_/Y _5114_/A _3876_/Y vssd1 vssd1 vccd1 vccd1 _3877_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2828_ _2826_/X _2717_/Y _2827_/X vssd1 vssd1 vccd1 vccd1 _2834_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__4360__A _4360_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5616_ _5692_/CLK _5616_/D vssd1 vssd1 vccd1 vccd1 _5616_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3176__A1 _5407_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5547_ _5641_/CLK _5547_/D vssd1 vssd1 vccd1 vccd1 _5547_/Q sky130_fd_sc_hd__dfxtp_1
X_2759_ _2916_/A _2864_/A _2759_/C _2864_/B vssd1 vssd1 vccd1 vccd1 _2852_/D sky130_fd_sc_hd__nand4_2
XANTENNA__5606__D _5606_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5478_ _5482_/CLK _5478_/D vssd1 vssd1 vccd1 vccd1 _5478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429_ _5264_/C vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3704__A _4057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5191__A _5200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3423__B _3433_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5341__D _5341_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4535__A _4535_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A2 _2927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A ksc_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4254__B _4265_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3939__B1 _3938_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4701__C _4716_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input74_A gpio_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5516__D _5516_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3614__A _3614_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2678__B1 _2677_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output230_A _3322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4419__A1 _2826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output328_A _3614_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5092__A1 _5081_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4445__A _4445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3992__A2_N _5673_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3800_ _3720_/X _3722_/X _3798_/X _3799_/X _3740_/X vssd1 vssd1 vccd1 vccd1 _3800_/Y
+ sky130_fd_sc_hd__o221ai_2
X_4780_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__C1 _3946_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3731_ _4099_/A vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3662_ _2771_/A _3998_/A _5590_/Q vssd1 vssd1 vccd1 vccd1 _3662_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__4611__C _5017_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3158__A1 _5404_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5401_ _5446_/CLK _5401_/D vssd1 vssd1 vccd1 vccd1 _5401_/Q sky130_fd_sc_hd__dfxtp_1
X_2613_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__buf_6
X_3593_ _4340_/B _5611_/Q _3600_/S vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5426__D _5426_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2905__A1 _2690_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5332_ _5737_/CLK _5332_/D vssd1 vssd1 vccd1 vccd1 _5332_/Q sky130_fd_sc_hd__dfxtp_1
X_2544_ _2544_/A _2544_/B _2583_/A _2581_/A vssd1 vssd1 vccd1 vccd1 _2640_/A sky130_fd_sc_hd__nand4_4
XFILLER_86_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _2667_/Y _5227_/A _2668_/Y vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__o21ai_1
XFILLER_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3524__A _3526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4214_ _4240_/A _4214_/B _4240_/C _4214_/D vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__and4_2
XFILLER_25_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2669__B1 _2668_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5194_ _5194_/A vssd1 vssd1 vccd1 vccd1 _5728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4145_ _4145_/A _4228_/B _4145_/C vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__and3_1
XFILLER_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3881__A2 _5774_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4058__C _4159_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4076_ _4076_/A vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5083__A1 _5075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3027_ _3027_/A _5444_/Q vssd1 vssd1 vccd1 vccd1 _3028_/A sky130_fd_sc_hd__and2_1
XANTENNA__4355__A _4355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4978_ _4978_/A _4997_/B _4997_/C vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__and3_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5240__D1 _5236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4594__B1 _4584_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3929_ _5777_/Q _3915_/X _3918_/X _3928_/Y vssd1 vssd1 vccd1 vccd1 _3930_/B sky130_fd_sc_hd__o22ai_4
XFILLER_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5186__A _5200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4090__A _4123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3149__A1 input42/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5336__D _5336_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4240__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3434__A _3434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4249__B _4249_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2695__D _2695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5522__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2992__B _5428_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5074__A1 _4889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3085__A0 _5143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__A _4265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5672__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__B1 _2831_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__C1 _4007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4585__B1 _4584_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4712__B _4731_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5096__A _5096_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__C1 _2691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4431__C _4431_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output180_A _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output278_A _3452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4888__A1 _3662_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3344__A _3344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5301__A2 _5268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4159__B _4159_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3863__A2 _3766_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5065__A1 _5662_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5065__B2 _5065_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4273__C1 _4272_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4901_ _4913_/A _4913_/B _4901_/C vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__or3_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2823__B1 _5380_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4903__A _4903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4832_ _5090_/A vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__buf_2
XFILLER_72_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3379__A1 _5503_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4763_ _4771_/A _4763_/B _4763_/C vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__or3_1
XFILLER_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4622__B _4622_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3519__A _3519_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__C1 _2696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3714_ _3994_/A vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__buf_4
X_4694_ _4699_/A _4714_/B _4694_/C vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__or3_1
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3645_ _4373_/A _5626_/Q _3645_/S vssd1 vssd1 vccd1 vccd1 _4984_/C sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4879__A1 _4163_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4879__B2 _4873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3576_ _4329_/A _5606_/Q _3597_/S vssd1 vssd1 vccd1 vccd1 _4934_/C sky130_fd_sc_hd__mux2_1
XFILLER_66_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3551__A1 _5599_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5315_ _5765_/CLK _5315_/D vssd1 vssd1 vccd1 vccd1 _5315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5545__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3254__A _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2796__C _2796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4170__A1_N _4139_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5172__C _5172_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5246_ _5752_/Q _5234_/X _2813_/Y _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5752_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__4069__B _4069_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3884__A2_N _5667_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3839__C1 _3838_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5177_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2657__A3 _2695_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3854__A2 _4128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5695__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4128_ _4128_/A vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_1_1_CLK_A clkbuf_1_1_1_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3067__A0 _4308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3899__A2_N _5668_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4059_ _4059_/A vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__buf_4
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3420__C _4739_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2814__B1 _2813_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4016__C1 _4015_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4532__B _4556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3429__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__A2 _3958_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input176_A spi_err_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A cpu_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4707__B _4707_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2805__B1 _5371_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4270__A2 _3830_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3862__B_N _3861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4723__A _4723_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5418__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output395_A _3166_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3339__A _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3230__A0 _4371_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5568__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3430_ _3430_/A vssd1 vssd1 vccd1 vccd1 _3430_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2897__B _2925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3361_ _3376_/A _3361_/B _4699_/C vssd1 vssd1 vccd1 vccd1 _3362_/A sky130_fd_sc_hd__and3_1
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5704__D _5704_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3074__A _3074_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5099_/X _5094_/X _5087_/X _5084_/X _4127_/B vssd1 vssd1 vccd1 vccd1 _5681_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3292_ _3292_/A _5538_/Q vssd1 vssd1 vccd1 vccd1 _3293_/A sky130_fd_sc_hd__and2_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _5779_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4089__A2 _4070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5031_ _5043_/A _5645_/Q _5039_/C _5043_/D vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__and4_1
XFILLER_100_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__B2 _3964_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5038__A1 _5648_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4617__B _4617_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5038__B2 _5034_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4246__C1 _4835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4261__A2 _4255_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815_ _4815_/A vssd1 vssd1 vccd1 vccd1 _5547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5795_ _5802_/CLK _5795_/D vssd1 vssd1 vccd1 vccd1 _5795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5167__C _5167_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4746_ _4746_/A vssd1 vssd1 vccd1 vccd1 _4765_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4677_ _4677_/A vssd1 vssd1 vccd1 vccd1 _5489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3628_ _3628_/A vssd1 vssd1 vccd1 vccd1 _3628_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2600__B _2600_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3559_ _3559_/A vssd1 vssd1 vccd1 vccd1 _3559_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5614__D _5614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput106 gpio_err_i vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__clkbuf_2
Xinput117 ksc_dat_i[17] vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput128 ksc_dat_i[27] vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput139 ksc_dat_i[8] vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5229_ _2836_/Y _5227_/X _2628_/C _5228_/X _4377_/X vssd1 vssd1 vccd1 vccd1 _5743_/D
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__4808__A _4821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3712__A _4075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _4543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A2 _4003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3159__A _3183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5710__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2998__A _2998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3593__S _3600_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3606__B _3620_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5524__D _5524_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__C1 _2787_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4718__A _4776_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3622__A _3622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4437__B _4437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output310_A _3476_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output408_A _3069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3451__A0 _4299_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4453__A _5228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2930_ _4415_/A _4415_/B _2780_/B _2787_/A _2787_/B vssd1 vssd1 vccd1 vccd1 _2937_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5268__B _5268_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2861_ _5697_/Q vssd1 vssd1 vccd1 vccd1 _2861_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4172__B _4172_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5390__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3069__A _3069_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4600_ _4600_/A vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3203__A0 _5191_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5580_ _5586_/CLK _5580_/D vssd1 vssd1 vccd1 vccd1 _5580_/Q sky130_fd_sc_hd__dfxtp_1
X_2792_ _2610_/A _5227_/A _2791_/Y _2540_/X vssd1 vssd1 vccd1 vccd1 _2792_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4531_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4556_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5284__A _5284_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4462_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__clkbuf_4
X_3413_ _3413_/A vssd1 vssd1 vccd1 vccd1 _3413_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5434__D _5434_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4393_ _4393_/A vssd1 vssd1 vccd1 vccd1 _5355_/D sky130_fd_sc_hd__clkbuf_1
X_3344_ _3344_/A vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__clkbuf_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 _2639_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3275_ _4396_/B _5531_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4628__A _4628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3532__A _3699_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5021_/A _5637_/Q _5017_/C _5021_/D vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__and4_1
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__A2 _3722_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5733__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4363__A _4363_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5178__B _5178_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5609__D _5609_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5778_ _5800_/CLK _5778_/D vssd1 vssd1 vccd1 vccd1 _5778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3745__A1 _5769_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4729_ _4749_/A _4739_/B _4729_/C vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__or3_1
XANTENNA__3745__B2 _3744_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5194__A _5194_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3707__A _4059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2611__A _2611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3426__B _3433_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__D _5344_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4170__B2 _4141_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2720__A2 _2594_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4538__A _4538_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3442__A _3445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input139_A ksc_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4063__B_N _4000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3984__A1 _3940_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5519__D _5519_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3617__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output260_A _3424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output358_A _3006_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4161__A1 _4161_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5606__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4448__A _5204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3352__A _3352_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3060_ _3163_/A vssd1 vssd1 vccd1 vccd1 _3230_/S sky130_fd_sc_hd__buf_4
XANTENNA__5110__B1 _5268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5756__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3672__B1 _5693_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4216__A2 _4449_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4183__A _4195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3962_ _3961_/X _3737_/X _5567_/Q vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4614__C _5017_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _5765_/CLK _5701_/D vssd1 vssd1 vccd1 vccd1 _5701_/Q sky130_fd_sc_hd__dfxtp_1
X_2913_ _3345_/A vssd1 vssd1 vccd1 vccd1 _3418_/A sky130_fd_sc_hd__buf_2
XANTENNA__5429__D _5429_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3893_ _4830_/B _3737_/X _5563_/Q vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4911__A _4911_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5632_ _5694_/CLK _5632_/D vssd1 vssd1 vccd1 vccd1 _5632_/Q sky130_fd_sc_hd__dfxtp_1
X_2844_ _5590_/Q _4115_/A _3678_/A vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__o21bai_4
XFILLER_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5563_ _5802_/CLK _5563_/D vssd1 vssd1 vccd1 vccd1 _5563_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2775_ _5802_/Q vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__buf_4
XANTENNA__3527__A _3527_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4514_ _4514_/A _4524_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__or3_1
XFILLER_69_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5494_ _5538_/CLK _5494_/D vssd1 vssd1 vccd1 vccd1 _5494_/Q sky130_fd_sc_hd__dfxtp_1
X_4445_ _4445_/A _5102_/A _4542_/A vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__and3_1
XANTENNA__4152__A1 _4147_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4376_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5264_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2702__A2 _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3327_ _3329_/A _5554_/Q vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__and2_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__A _4358_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__B1 _5097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3258_ _3407_/A vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3189_ _3210_/A _3194_/B _4517_/A vssd1 vssd1 vccd1 vccd1 _3190_/A sky130_fd_sc_hd__and3_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3663__B1 _3678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4207__A2 _4115_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5189__A _5189_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3415__A0 _4353_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2606__A _2621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4524__C _4524_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2769__A2 _2879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5339__D _5339_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4243__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__A _4821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3718__A1 _3718_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3437__A _3437_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5629__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2698__D _2831_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5779__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5802__D _5802_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4268__A _5587_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3172__A _3172_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__A0 _4301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__A _4240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4851__C1 _4843_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__A _5099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4603__C1 _4598_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4731__A _4731_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _5695_/Q vssd1 vssd1 vccd1 vccd1 _2560_/Y sky130_fd_sc_hd__clkinv_2
Xoutput207 _3897_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput218 _3298_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput229 _3320_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[26] sky130_fd_sc_hd__buf_2
XFILLER_86_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4134__A1 _3997_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4134__B2 _4133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4230_ _5584_/Q vssd1 vssd1 vccd1 vccd1 _4230_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4161_ _4161_/A1 _4449_/A _3994_/A _4160_/Y vssd1 vssd1 vccd1 vccd1 _4654_/B sky130_fd_sc_hd__a31oi_4
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5712__D _5712_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3082__A _3082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3893__B1 _5563_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3112_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4092_ _4092_/A vssd1 vssd1 vccd1 vccd1 _4092_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5095__C1 _4094_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3043_ _3043_/A vssd1 vssd1 vccd1 vccd1 _3043_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3645__A0 _4373_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4906__A _4906_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3810__A _4171_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4994_ _5156_/A vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__buf_8
XANTENNA__3948__A1 _5778_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3948__B2 _3947_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3945_ _3940_/X _3825_/X _3826_/X _3944_/Y vssd1 vssd1 vccd1 vccd1 _3945_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4063__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4641__A _4645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2620__A1 _5359_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3876_ _4628_/A _3857_/X _5099_/A _3875_/Y vssd1 vssd1 vccd1 vccd1 _3876_/Y sky130_fd_sc_hd__o211ai_1
X_5615_ _5692_/CLK _5615_/D vssd1 vssd1 vccd1 vccd1 _5615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ _5759_/Q _2683_/X _2658_/Y _2574_/X vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4360__B _4381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3257__A _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5546_ _5555_/CLK _5546_/D vssd1 vssd1 vccd1 vccd1 _5546_/Q sky130_fd_sc_hd__dfxtp_1
X_2758_ _5364_/Q _2611_/A _2757_/Y vssd1 vssd1 vccd1 vccd1 _2916_/A sky130_fd_sc_hd__o21ai_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5477_ _5798_/CLK _5477_/D vssd1 vssd1 vccd1 vccd1 _5477_/Q sky130_fd_sc_hd__dfxtp_1
X_2689_ _2682_/Y _2565_/X _2688_/Y vssd1 vssd1 vccd1 vccd1 _2689_/Y sky130_fd_sc_hd__o21ai_2
X_4428_ _4428_/A vssd1 vssd1 vccd1 vccd1 _5373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5191__B _5191_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5622__D _5622_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4359_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3884__B1 _3883_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3423__C _4741_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5086__C1 _5064_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3636__A0 _4366_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3720__A _4147_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__C _4254_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _5462_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4061__B1 _4060_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4551__A _4551_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5451__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3167__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input67_A cpu_sel_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5532__D _5532_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2678__A1 _5266_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3875__B1 _3874_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4419__A2 _2717_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5077__C1 _3900_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2945__S _3233_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4726__A _4726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output223_A _3307_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3630__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4824__C1 _4823_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5092__A2 _5078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4445__B _5102_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__B1 _4051_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4461__A _4461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3730_ _3980_/A vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ _3980_/A _4082_/A _4083_/A _2800_/A vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__o31a_2
XANTENNA__5707__D _5707_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3077__A _3250_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4611__D _4614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5400_ _5731_/CLK _5400_/D vssd1 vssd1 vccd1 vccd1 _5400_/Q sky130_fd_sc_hd__dfxtp_1
X_2612_ _2605_/Y _2606_/X _2611_/Y vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__o21ai_2
X_3592_ _3592_/A vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2905__A2 _5195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5331_ _5741_/CLK _5331_/D vssd1 vssd1 vccd1 vccd1 _5331_/Q sky130_fd_sc_hd__dfxtp_1
X_2543_ _2543_/A vssd1 vssd1 vccd1 vccd1 _2544_/B sky130_fd_sc_hd__buf_2
XANTENNA__3805__A _5068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5262_ _2709_/Y _5261_/X _4565_/X _4400_/X vssd1 vssd1 vccd1 vccd1 _5765_/D sky130_fd_sc_hd__a211o_1
XFILLER_69_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3524__B _5656_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4213_ _3806_/X _5687_/Q _4212_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _4214_/B sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__2669__A1 _2667_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5442__D _5442_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5193_ _5193_/A _5202_/B _5208_/C vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__and3_1
XFILLER_69_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4144_ _4075_/X _4076_/X _4144_/C _4201_/D vssd1 vssd1 vccd1 vccd1 _4145_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__4213__A2_N _5687_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5324__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4058__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4636__A _4638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4075_ _4075_/A vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3540__A _3540_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5083__A2 _4890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3026_ _3026_/A vssd1 vssd1 vccd1 vccd1 _3026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4355__B _4355_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5474__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4977_ _4977_/A vssd1 vssd1 vccd1 vccd1 _5622_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5240__C1 _5235_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4594__A1 _5440_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4371__A _4396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4594__B2 _4590_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3928_ _3887_/X _4636_/B _3927_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _3928_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_36_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5186__B _5191_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4090__B _5295_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5617__D _5617_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3859_ _5561_/Q vssd1 vssd1 vccd1 vccd1 _3859_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529_ _5531_/CLK _5529_/D vssd1 vssd1 vccd1 vccd1 _5529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3715__A _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5352__D _5352_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3609__A0 _4349_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4546__A _4546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4806__C1 _4805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5074__A2 _5060_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input121_A ksc_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3085__A1 _5322_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4282__B1 _4281_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__B _4265_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2832__A1 _5754_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4034__B1 _4033_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4585__A1 _5436_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4585__B2 _4564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4712__C _4716_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__B1 _2595_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5527__D _5527_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4888__A2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3625__A _3625_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5298__C1 _5278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5347__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output340_A _3548_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4159__C _4159_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4456__A _4891_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5497__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5065__A2 _4988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4273__B1 _4267_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _4968_/A vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2823__A1 _2809_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4831_ _4831_/A vssd1 vssd1 vccd1 vccd1 _5556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4903__B _4915_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5287__A _5287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _5523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2704__A _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2587__B1 _2585_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3713_ _4265_/C vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5437__D _5437_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4693_ _4776_/B vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3644_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4879__A2 _4164_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3575_ _3575_/A vssd1 vssd1 vccd1 vccd1 _3575_/X sky130_fd_sc_hd__clkbuf_1
X_5314_ _5741_/CLK _5314_/D vssd1 vssd1 vccd1 vccd1 _5314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5244_/X _2648_/Y _4891_/X _5238_/X vssd1 vssd1 vccd1 vccd1 _5751_/D sky130_fd_sc_hd__a211o_1
XFILLER_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3839__B1 _3826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5176_ _5176_/A _5191_/B _5176_/C vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__or3_1
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4127_ _4127_/A _4127_/B _4159_/C _4214_/D vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__and4_2
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4366__A _4366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3067__A1 _5389_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4058_ _4127_/A _4058_/B _4159_/C _4214_/D vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__and4_2
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4264__B1 _3846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3009_ _3009_/A vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2814__A1 _5752_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4016__B1 _5099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5197__A _5197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2614__A _2614_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4532__C _4536_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3429__B _3433_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3775__C1 _3774_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5347__D _5347_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3445__A _3445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input169_A spi_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput390 _3135_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_43_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4707__C _4716_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4255__B1 _4254_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2805__A1 _2569_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3339__B _4761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output290_A _3501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3230__A1 _5417_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output388_A _3124_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3355__A _3355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2897__C _2911_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3360_ _4320_/A _5498_/Q _3441_/S vssd1 vssd1 vccd1 vccd1 _4699_/C sky130_fd_sc_hd__mux2_1
XFILLER_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3291_/X sky130_fd_sc_hd__clkbuf_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5286__A2 _5269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5030_ _5644_/Q _5010_/X _5029_/X _5011_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5644_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5720__D _5720_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5038__A2 _5033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4617__C _4796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4246__B1 _4244_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4914__A _4914_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _4821_/A _5547_/Q _4817_/C vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__and3_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5794_ _5798_/CLK _5794_/D vssd1 vssd1 vccd1 vccd1 _5794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _5516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5512__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4676_ _4676_/A _4681_/B _4690_/C vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__and3_1
XANTENNA__2980__A0 _5221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3627_ _3630_/A _3637_/B _4969_/C vssd1 vssd1 vccd1 vccd1 _3628_/A sky130_fd_sc_hd__and3_1
XFILLER_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3558_ _3558_/A _3565_/B _4924_/A vssd1 vssd1 vccd1 vccd1 _3559_/A sky130_fd_sc_hd__and3_1
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5662__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2600__C _2600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2732__B1 _4417_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3489_ _3493_/A _5640_/Q vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__and2_1
XFILLER_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput107 gpio_rty_i vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput118 ksc_dat_i[18] vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5228_ _5228_/A vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__buf_2
Xinput129 ksc_dat_i[28] vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4808__B _5543_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3712__B _4076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2609__A input5/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5159_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5630__D _5630_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3204__S _3204_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3159__B _3165_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2971__A0 _4388_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3606__C _4955_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__B1 _2782_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3903__A _4283_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5540__D _5540_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4437__C _4437_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output303_A _3527_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4734__A _4734_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3451__A1 _5489_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5535__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2860_ _2751_/Y _2574_/X _2850_/D vssd1 vssd1 vccd1 vccd1 _2916_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__5268__C _5268_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4172__C _4252_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3203__A1 _5342_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2791_ _5261_/B _2708_/X _5747_/Q vssd1 vssd1 vccd1 vccd1 _2791_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _4530_/A vssd1 vssd1 vccd1 vccd1 _5414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5685__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5284__B _5284_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2962__B1 _4548_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4461_ _4461_/A vssd1 vssd1 vccd1 vccd1 _5388_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5715__D _5715_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3412_ _3412_/A _3416_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _3413_/A sky130_fd_sc_hd__and3_1
X_4392_ _4396_/A _4392_/B vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__and2_1
XANTENNA__2714__B1 _4431_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3911__C1 _3910_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3343_ _3357_/A _4761_/A _4686_/A vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__and3_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__A _4913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A2 _5227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3813__A _4059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3267_/X _3268_/X _4776_/C vssd1 vssd1 vccd1 vccd1 _3274_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5013_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__buf_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__D _5450_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4219__B1 _5583_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4644__A _4651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5178__C _5184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5777_ _5800_/CLK _5777_/D vssd1 vssd1 vccd1 vccd1 _5777_/Q sky130_fd_sc_hd__dfxtp_1
X_2989_ _4396_/B _5427_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__mux2_1
X_4728_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3745__A2 _3690_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5625__D _5625_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2611__B _2611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4659_ _5480_/Q _4652_/X _4228_/X _4621_/A vssd1 vssd1 vccd1 vccd1 _5480_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3426__C _4744_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3723__A _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5408__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4538__B _4550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3442__B _3445_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5360__D _5360_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4257__C _4257_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5558__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4554__A _4674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3984__A2 _3825_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input97_A gpio_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3197__A0 _5726_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3617__B _3620_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5535__D _5535_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3109__S _3132_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2948__S _3234_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4161__A2 _4449_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output253_A _3402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4729__A _4749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5110__A1 _5096_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output420_A _3249_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3121__A0 _5157_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3672__A1 _5058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4464__A _4464_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4216__A3 _3994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4183__B _5302_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _3961_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__D _4614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5700_ _5766_/CLK _5700_/D vssd1 vssd1 vccd1 vccd1 _5700_/Q sky130_fd_sc_hd__dfxtp_1
X_2912_ _2900_/Y _2910_/Y _2911_/Y vssd1 vssd1 vccd1 vccd1 _3345_/A sky130_fd_sc_hd__o21ai_4
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3892_ _3277_/A _3723_/X _3725_/X _3891_/X vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__o211a_1
X_5631_ _5641_/CLK _5631_/D vssd1 vssd1 vccd1 vccd1 _5631_/Q sky130_fd_sc_hd__dfxtp_1
X_2843_ _5696_/Q _3957_/A _5802_/Q vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__4911__B _4915_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3188__A0 _4353_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5295__A _5295_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3808__A _4141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5562_ _5589_/CLK _5562_/D vssd1 vssd1 vccd1 vccd1 _5562_/Q sky130_fd_sc_hd__dfxtp_1
X_2774_ _4830_/A vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__buf_2
XFILLER_34_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4513_ _4513_/A vssd1 vssd1 vccd1 vccd1 _5407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5445__D _5445_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5493_ _5538_/CLK _5493_/D vssd1 vssd1 vccd1 vccd1 _5493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__buf_4
XFILLER_67_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4152__A2 _4046_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4639__A _4652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3360__A0 _4320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3326_/A vssd1 vssd1 vccd1 vccd1 _3326_/X sky130_fd_sc_hd__clkbuf_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5101__A1 _5096_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3257_ _3403_/A vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__clkbuf_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5700__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3188_ _4353_/B _5409_/Q _3209_/S vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3663__A1 _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3663__B2 _3662_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4162__A_N _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4374__A _4374_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5189__B _5202_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3415__A1 _5513_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2769__A3 _2909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4821__B _5551_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2622__A _2622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3718__A2 _4528_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5355__D _5355_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4549__A _4549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input151_A spi_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4030__B_N _4000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5380__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__A1 _5594_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A cpu_adr_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4851__B1 _4832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3900__B _3900_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2862__C1 _2859_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4603__B1 _4584_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4731__B _4731_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3628__A _3628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output370_A _3031_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3590__A0 _4338_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput208 _3914_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput219 _3300_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4134__A2 _4062_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4459__A _4459_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5723__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3363__A _3418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3342__A0 _4308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4160_ _4027_/X _4095_/X _5475_/Q vssd1 vssd1 vccd1 vccd1 _4160_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__3893__A1 _4830_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3111_ _3123_/A _3134_/B _4483_/C vssd1 vssd1 vccd1 vccd1 _3112_/A sky130_fd_sc_hd__and3_1
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _4091_/X sky130_fd_sc_hd__buf_4
XANTENNA__5095__B1 _5084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3042_ _3042_/A _5451_/Q vssd1 vssd1 vccd1 vccd1 _3043_/A sky130_fd_sc_hd__and2_1
XANTENNA__3645__A1 _5626_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2707__A _2707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4993_ _4993_/A vssd1 vssd1 vccd1 vccd1 _5629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4922__A _4947_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3948__A2 _3804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3944_ _3941_/Y _3906_/X _3943_/Y vssd1 vssd1 vccd1 vccd1 _3944_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _3872_/Y _4743_/A _3874_/Y vssd1 vssd1 vccd1 vccd1 _3875_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2620__A2 _2613_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3538__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5614_ _5692_/CLK _5614_/D vssd1 vssd1 vccd1 vccd1 _5614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2826_ _2806_/X _5266_/A _5368_/Q vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5545_ _5641_/CLK _5545_/D vssd1 vssd1 vccd1 vccd1 _5545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2757_ _2592_/Y _2790_/A _2595_/Y _2704_/A _2806_/A vssd1 vssd1 vccd1 vccd1 _2757_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_69_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5476_ _5482_/CLK _5476_/D vssd1 vssd1 vccd1 vccd1 _5476_/Q sky130_fd_sc_hd__dfxtp_1
X_2688_ _5758_/Q _2683_/X _2687_/Y _2574_/X vssd1 vssd1 vccd1 vccd1 _2688_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4427_ _4431_/A _4427_/B _4427_/C vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__and3_1
XANTENNA__4369__A _4369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5191__C _5191_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _5341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A cpu_adr_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3884__B2 _3700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3309_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3309_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4295_/C _4567_/A _4407_/A _4289_/D vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__and4b_4
XANTENNA__5086__B1 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3636__A1 _5623_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2617__A _2652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4832__A _5090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3939__A2 _3815_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4061__A1 _4061_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5746__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3183__A _3183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2678__A2 _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3875__A1 _3872_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5077__B1 _5076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4726__B _4731_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4824__B1 _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3630__B _3637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5092__A3 _5087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output216_A _3293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3122__S _3146_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4445__C _4542_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2961__S _3240_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4742__A _4742_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__A1 _4042_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3358__A _3358_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3660_ _3660_/A vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2611_ _2611_/A _2611_/B _2611_/C vssd1 vssd1 vccd1 vccd1 _2611_/Y sky130_fd_sc_hd__nand3_1
X_3591_ _3594_/A _3601_/B _4945_/C vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__and3_1
XFILLER_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5330_ _5741_/CLK _5330_/D vssd1 vssd1 vccd1 vccd1 _5330_/Q sky130_fd_sc_hd__dfxtp_1
X_2542_ _5768_/Q vssd1 vssd1 vccd1 vccd1 _2544_/A sky130_fd_sc_hd__inv_2
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A _5261_/B _5261_/C _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__or4_1
XANTENNA__5723__D _5723_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3093__A _3093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__inv_2
X_5192_ _5192_/A vssd1 vssd1 vccd1 vccd1 _5727_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2669__A2 _2640_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _4252_/A _4143_/B _4143_/C _4172_/D vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__and4_4
XANTENNA__4917__A _4917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3821__A _4283_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4074_ _4074_/A vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4636__B _4636_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3540__B _3547_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3027_/A _5443_/Q vssd1 vssd1 vccd1 vccd1 _3026_/A sky130_fd_sc_hd__and2_1
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5083__A3 _5070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5619__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4652__A _4652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4976_ _4990_/A _4990_/B _4976_/C vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__or3_1
XANTENNA__5240__B1 _2585_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4594__A2 _4589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3927_ _3720_/X _3890_/X _3925_/X _3926_/X _3740_/X vssd1 vssd1 vccd1 vccd1 _3927_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4371__B _4371_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5769__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3268__A _4295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5186__C _5186_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3858_ _4005_/A vssd1 vssd1 vccd1 vccd1 _4835_/A sky130_fd_sc_hd__clkbuf_4
X_2809_ _2809_/A vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__clkbuf_4
X_3789_ _3695_/X _5663_/Q _3788_/Y _3700_/X vssd1 vssd1 vccd1 vccd1 _3792_/B sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__3554__A0 _4316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2900__A _5523_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5528_ _5635_/CLK _5528_/D vssd1 vssd1 vccd1 vccd1 _5528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2762__D1 _2806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4099__A _4099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5459_ _5741_/CLK _5459_/D vssd1 vssd1 vccd1 vccd1 _5459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5633__D _5633_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3207__S _3228_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3731__A _4099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3609__A1 _5615_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__B1 _4798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5074__A3 _5066_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4282__A1 _4276_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__C _4265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input114_A ksc_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__A2 _2683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4562__A _4562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__A1 _3887_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4585__A2 _4563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3178__A _3178_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__A1 _2707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3906__A _4692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4888__A3 _4847_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5543__D _5543_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5298__B1 _4127_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4159__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4737__A _4737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output333_A _3631_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3641__A _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4456__B _4473_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__D1 _4117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4273__A1 _5111_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2823__A2 _2750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4472__A _4472_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _4830_/A _4830_/B _4988_/C vssd1 vssd1 vccd1 vccd1 _4831_/A sky130_fd_sc_hd__and3_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4903__C _4915_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4761_ _4761_/A _4778_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__and3_1
XFILLER_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5718__D _5718_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3088__A _3088_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__A1 _5748_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3712_ _4075_/A _4076_/A _4253_/D vssd1 vssd1 vccd1 vccd1 _4265_/C sky130_fd_sc_hd__nor3b_2
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4692_ _4692_/A vssd1 vssd1 vccd1 vccd1 _4776_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3643_ _3646_/A _4988_/B _4982_/A vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__and3_1
XANTENNA__3816__A _3849_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3574_ _3577_/A _3584_/B _4932_/A vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__and3_1
X_5313_ _5765_/CLK _5313_/D vssd1 vssd1 vccd1 vccd1 _5313_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5453__D _5453_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5244_ _2813_/C _2831_/D _2831_/B _5751_/Q vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3839__A1 _3824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5175_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5720_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4647__A _4651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5441__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4126_ _3989_/X _5681_/Q _4125_/Y _3991_/X vssd1 vssd1 vccd1 vccd1 _4127_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_99_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4366__B _4366_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A vssd1 vssd1 vccd1 vccd1 _4214_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4264__A1 _5691_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4264__B2 _4264_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3008_ _3016_/A _5435_/Q vssd1 vssd1 vccd1 vccd1 _3009_/A sky130_fd_sc_hd__and2_1
XANTENNA__2814__A2 _2683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5591__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4382__A _4382_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4016__A1 _4628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4959_ _4963_/A _4963_/B _4959_/C vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__or3_1
XFILLER_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5628__D _5628_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__B1 _5099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3429__C _4747_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3959__B_N _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3726__A _4082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__A _4405_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3445__B _3445_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5363__D _5363_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput380 _2982_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[5] sky130_fd_sc_hd__buf_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3955__B1_N _5463_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput391 _3142_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4557__A _4557_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4255__A1 _5482_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2805__A2 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4292__A _4299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3400__S _3400_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__D _5538_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3339__C _4683_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output283_A _3486_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5314__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2540__A _2691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4191__B1 _4190_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5464__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3290_ _3292_/A _5537_/Q vssd1 vssd1 vccd1 vccd1 _3291_/A sky130_fd_sc_hd__and2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4467__A _5270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3371__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4246__A1 _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4246__B2 _4245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2715__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4813_ _5546_/Q _4803_/X _4798_/X _4804_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5546_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5448__D _5448_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5793_ _5802_/CLK _5793_/D vssd1 vssd1 vccd1 vccd1 _5793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4930__A _4938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4744_ _4749_/A _4763_/B _4744_/C vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__or3_1
XFILLER_33_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4675_ _4675_/A vssd1 vssd1 vccd1 vccd1 _5488_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2980__A1 _5355_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3626_ _4360_/A _5620_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _4969_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2717__D1 _2672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4182__B1 _4172_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3557_ _4318_/B _5601_/Q _3564_/S vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2732__A1 _5367_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4269__A_N _3860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__clkbuf_1
Xinput108 ksc_ack_i vssd1 vssd1 vccd1 vccd1 _3670_/A1 sky130_fd_sc_hd__buf_2
X_5227_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__clkbuf_4
Xinput119 ksc_dat_i[19] vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4377__A _5264_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3281__A _3281_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4808__C _4817_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5158_ _5158_/A vssd1 vssd1 vccd1 vccd1 _5713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4109_ _4109_/A _4109_/B _4143_/C _4172_/D vssd1 vssd1 vccd1 vccd1 _4109_/X sky130_fd_sc_hd__and4_4
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _5089_/A vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2625__A _2684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3996__B1 _3995_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3220__S _3230_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5001__A _5183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5358__D _5358_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5337__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3159__C _4503_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4840__A _5268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3456__A _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2971__A1 _5423_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5487__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__A1 _4439_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A cpu_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3903__B _4079_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4287__A _4287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2535__A _5767_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5268__D _5268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4172__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4750__A _4750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2790_ _2790_/A vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3366__A _3366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2962__A1 _2876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4460_ _4891_/A _4473_/B _4460_/C vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_16_CLK clkbuf_opt_3_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5659_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3411_ _4351_/A _5512_/Q _3432_/S vssd1 vssd1 vccd1 vccd1 _4733_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4164__B1 _5579_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4391_ _4391_/A vssd1 vssd1 vccd1 vccd1 _5354_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2714__A1 _5375_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3342_ _4308_/B _5493_/Q _3364_/S vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3911__B1 _3826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4909__B _4913_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__C1 _3674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3273_ _4394_/A _5530_/Q _3453_/S vssd1 vssd1 vccd1 vccd1 _4776_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4197__A _4197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5731__D _5731_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5012_ _5636_/Q _5010_/X _5806_/A _5011_/X _4823_/X vssd1 vssd1 vccd1 vccd1 _5636_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4925__A _4925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4219__A1 _3735_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4644__B _4644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4660__A _4660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5776_ _5800_/CLK _5776_/D vssd1 vssd1 vccd1 vccd1 _5776_/Q sky130_fd_sc_hd__dfxtp_1
X_2988_ _5225_/A _5357_/Q _3229_/S vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__mux2_8
XFILLER_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4727_ _4727_/A vssd1 vssd1 vccd1 vccd1 _5509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4658_ _4660_/A _4658_/B vssd1 vssd1 vccd1 vccd1 _5479_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2611__C _2611_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput90 gpio_dat_i[24] vssd1 vssd1 vccd1 vccd1 _4189_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4155__B1 _4143_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3609_ _4349_/B _5615_/Q _3636_/S vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__mux2_1
X_4589_ _4600_/A vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5104__C1 _4172_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5641__D _5641_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3215__S _3235_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4538__C _4538_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3442__C _4756_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4257__D _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4835__A _4835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4554__B _4558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2641__B1 _5763_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4570__A _4570_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3197__A1 input51/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3617__C _4961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4146__B1 _4145_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3914__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__A3 _3994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4729__B _4739_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5551__D _5551_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output246_A _3377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5110__A2 _4837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3121__A1 _5328_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5502__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output413_A _3088_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4745__A _4745_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3672__A2 _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_5_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5737_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4464__B _4475_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3960_ _3922_/X _3958_/X _3725_/X _3959_/X vssd1 vssd1 vccd1 vccd1 _3960_/X sky130_fd_sc_hd__o211a_2
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5652__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _2886_/Y _2911_/B _2925_/B _2925_/A vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__nand4b_2
X_3891_ _3727_/X _3729_/X _3891_/C _3978_/A vssd1 vssd1 vccd1 vccd1 _3891_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4480__A _5228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2842_ _2842_/A _2842_/B _2842_/C vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__nor3_4
X_5630_ _5694_/CLK _5630_/D vssd1 vssd1 vccd1 vccd1 _5630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4911__C _4915_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3188__A1 _5409_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5295__B _5297_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2773_ _3331_/A vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__clkbuf_4
X_5561_ _5589_/CLK _5561_/D vssd1 vssd1 vccd1 vccd1 _5561_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5726__D _5726_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4512_ _4512_/A _4526_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__and3_1
XFILLER_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5492_ _5538_/CLK _5492_/D vssd1 vssd1 vccd1 vccd1 _5492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4443_ _2700_/X _2676_/X _4402_/X vssd1 vssd1 vccd1 vccd1 _5382_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__3824__A _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4374_ _4374_/A vssd1 vssd1 vccd1 vccd1 _5348_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3360__A1 _5498_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3325_ _3325_/A _5553_/Q vssd1 vssd1 vccd1 vccd1 _3326_/A sky130_fd_sc_hd__and2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5461__D _5461_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3256_ _2895_/X _2899_/X _4763_/C vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__o21a_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__A2 _5089_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3187_ _5184_/A _5339_/Q _3219_/S vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__mux2_8
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3663__A2 _3755_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2871__B1 _2870_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5189__C _5208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2769__A4 _2768_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4390__A _4390_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2903__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4821__C _4988_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5636__D _5636_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5759_ _5765_/CLK _5759_/D vssd1 vssd1 vccd1 vccd1 _5759_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3718__A3 _3714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3734__A _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5525__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5371__D _5371_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input144_A spi_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4565__A _4891_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4851__A1 _3892_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5675__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4851__B2 _4833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3900__C _4240_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2862__B1 _2861_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4064__C1 _4063_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4603__A1 _5444_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4603__B2 _4590_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2813__A _2813_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4198__A1_N _4139_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4731__C _4741_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5546__D _5546_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output196_A _4211_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3590__A1 _5610_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4119__B1 _4118_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput209 _3930_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[8] sky130_fd_sc_hd__buf_2
XANTENNA_output363_A _3017_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3644__A _3644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3342__A1 _5493_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _4324_/A _5396_/Q _3146_/S vssd1 vssd1 vccd1 vccd1 _4483_/C sky130_fd_sc_hd__mux2_1
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3893__A2 _3737_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _4123_/A _5295_/A vssd1 vssd1 vccd1 vccd1 _4090_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5095__A1 _5081_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3041_ _3041_/A vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4475__A _4475_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4992_ _4992_/A _4997_/B _4997_/C vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__and3_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5252__D1 _5236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3943_ _3829_/X _3830_/X _3831_/X _3942_/X _3908_/X vssd1 vssd1 vccd1 vccd1 _3943_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3819__A _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3874_ _3763_/X _3766_/X _3768_/X _3873_/X _3331_/A vssd1 vssd1 vccd1 vccd1 _3874_/Y
+ sky130_fd_sc_hd__o2111ai_1
X_5613_ _5692_/CLK _5613_/D vssd1 vssd1 vccd1 vccd1 _5613_/Q sky130_fd_sc_hd__dfxtp_1
X_2825_ _2823_/Y _2745_/Y _4431_/C _4431_/B vssd1 vssd1 vccd1 vccd1 _2908_/C sky130_fd_sc_hd__a22oi_4
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5456__D _5456_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5544_ _5555_/CLK _5544_/D vssd1 vssd1 vccd1 vccd1 _5544_/Q sky130_fd_sc_hd__dfxtp_1
X_2756_ _2752_/Y _2552_/Y _2755_/Y vssd1 vssd1 vccd1 vccd1 _2909_/C sky130_fd_sc_hd__a21oi_4
XFILLER_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5307__C1 _5278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5548__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2687_ _2734_/C _2831_/B _2813_/C _2831_/D vssd1 vssd1 vccd1 vccd1 _2687_/Y sky130_fd_sc_hd__nand4b_2
X_5475_ _5482_/CLK _5475_/D vssd1 vssd1 vccd1 vccd1 _5475_/Q sky130_fd_sc_hd__dfxtp_1
X_4426_ _4426_/A vssd1 vssd1 vccd1 vccd1 _5372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4357_ _4366_/A _4357_/B vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__and2_1
XFILLER_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5698__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3308_ _3314_/A _5545_/Q vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__and2_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ input1/X vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5086__A1 _5674_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5086__B2 _5086_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3239_ _5120_/A _5313_/Q _4375_/A vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4385__A _4385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4061__A2 _3954_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3729__A _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5366__D _5366_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3183__B _3194_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3875__A2 _4743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5077__A1 _5075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4295__A _4466_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4824__A1 _5552_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4726__C _4741_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4824__B2 _4804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3630__C _4974_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2835__B1 _5358_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output209_A _3930_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__A2 _4045_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2543__A _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3260__B1 _4765_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2610_ _2610_/A _2848_/B _2848_/C _2848_/D vssd1 vssd1 vccd1 vccd1 _2611_/C sky130_fd_sc_hd__nand4_2
X_3590_ _4338_/A _5610_/Q _3597_/S vssd1 vssd1 vccd1 vccd1 _4945_/C sky130_fd_sc_hd__mux2_1
XFILLER_70_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2541_ input3/X vssd1 vssd1 vccd1 vccd1 _2848_/A sky130_fd_sc_hd__inv_2
XFILLER_66_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3374__A _3374_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5260_ _5764_/Q _5234_/A _2698_/Y _5228_/X _4377_/X vssd1 vssd1 vccd1 vccd1 _5764_/D
+ sky130_fd_sc_hd__o2111a_1
X_4211_ _4263_/A _5304_/A vssd1 vssd1 vccd1 vccd1 _4211_/Y sky130_fd_sc_hd__nor2_8
XFILLER_9_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3789__A2_N _5663_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5191_ _5200_/A _5191_/B _5191_/C vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__or3_1
X_4142_ _4139_/X _5682_/Q _4140_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _4143_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3079__A0 _5141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3821__B _4283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4073_ _4109_/A _4073_/B _4143_/C _4172_/D vssd1 vssd1 vccd1 vccd1 _4073_/X sky130_fd_sc_hd__and4_4
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3024_ _3024_/A vssd1 vssd1 vccd1 vccd1 _3024_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3540__C _4909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2826__B1 _5368_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4933__A _4933_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _4975_/A vssd1 vssd1 vccd1 vccd1 _5621_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5240__A1 _5748_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3549__A _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3251__A0 _5128_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3926_ _4830_/B _3737_/X _5565_/Q vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5370__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3857_ _3857_/A vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2808_ _4423_/C _4423_/B _4441_/C _4441_/B vssd1 vssd1 vccd1 vccd1 _2902_/D sky130_fd_sc_hd__a22oi_4
X_3788_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3788_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3554__A1 _5600_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5527_ _5531_/CLK _5527_/D vssd1 vssd1 vccd1 vccd1 _5527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2739_ _2621_/X _2696_/B _2696_/C _4421_/A vssd1 vssd1 vccd1 vccd1 _2780_/D sky130_fd_sc_hd__a31oi_4
XANTENNA__3284__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2762__C1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5458_ _5798_/CLK _5458_/D vssd1 vssd1 vccd1 vccd1 _5458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4409_ _4567_/A vssd1 vssd1 vccd1 vccd1 _5228_/A sky130_fd_sc_hd__buf_6
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5389_ _5435_/CLK _5389_/D vssd1 vssd1 vccd1 vccd1 _5389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2628__A _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3223__S _3223_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__A1 _5542_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5004__A _5004_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4806__B2 _4804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2817__B1 _5378_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4282__A2 _3848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__D _4265_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4843__A _5235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A gpio_rty_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4034__A2 _4644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3459__A _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5713__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3242__A0 _5699_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__A2 _2592_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input72_A cpu_we_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3194__A _3210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5298__A1 _5789_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5298__B2 _4135_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__A _4098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4737__B _4756_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2538__A _2573_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output326_A _3541_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3133__S _3146_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4258__C1 _4257_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4456__C _4456_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2808__B1 _4441_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4273__A2 _3848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4753__A _4917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4043__B_N _3818_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5393__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3369__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3233__A0 _5733_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4760_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__C1 _4402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2587__A2 _2577_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3711_ _3711_/A vssd1 vssd1 vccd1 vccd1 _4253_/D sky130_fd_sc_hd__clkbuf_2
X_4691_ _4691_/A vssd1 vssd1 vccd1 vccd1 _5495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3642_ _4371_/B _5625_/Q _3642_/S vssd1 vssd1 vccd1 vccd1 _4982_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3573_ _4327_/B _5605_/Q _3600_/S vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5734__D _5734_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5312_ _5268_/B _5096_/A _5114_/X _5102_/X _5268_/C vssd1 vssd1 vccd1 vccd1 _5802_/D
+ sky130_fd_sc_hd__o311a_1
X_5243_ _2600_/B _2600_/C _5242_/Y vssd1 vssd1 vccd1 vccd1 _5750_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__4928__A _4928_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3832__A _4082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3839__A2 _3825_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5174_ _5174_/A _5178_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__and3_1
XFILLER_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4647__B _4647_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4125_ _4125_/A vssd1 vssd1 vccd1 vccd1 _4125_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4048__A_N _3832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _3989_/X _5677_/Q _4055_/Y _3991_/X vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4264__A2 _4986_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3007_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3016_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5736__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3472__B1 _4999_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4016__A2 _3857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3279__A _3281_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3224__A0 _5200_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ _4958_/A vssd1 vssd1 vccd1 vccd1 _5615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3775__A1 _4628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3909_ _3829_/X _3830_/X _3831_/X _3907_/X _3908_/X vssd1 vssd1 vccd1 vccd1 _3909_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_32_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4889_ _5081_/A vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5644__D _5644_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__B _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_7_CLK_A clkbuf_leaf_7_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3218__S _3228_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3445__C _4758_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4838__A _5270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput370 _3031_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput381 _2986_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__3742__A _3742_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput392 _3148_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4255__A2 _4489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4573__A _4592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3463__A0 _4386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__B _4292_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3189__A _3210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__A0 _4364_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output276_A _3448_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5554__D _5554_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3128__S _3151_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4191__A1 _4188_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5609__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__A _4748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5759__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4246__A2 _3857_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4483__A _4487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3454__B1 _4679_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5729__D _5729_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3099__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4812_ _4812_/A vssd1 vssd1 vccd1 vccd1 _5545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5792_ _5798_/CLK _5792_/D vssd1 vssd1 vccd1 vccd1 _5792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743_ _4743_/A vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4930__B _4938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3827__A _5560_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4674_ _4674_/A _4688_/B _4674_/C vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__or3_1
X_3625_ _3625_/A vssd1 vssd1 vccd1 vccd1 _3625_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5464__D _5464_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2717__C1 _2699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4182__A1 _5792_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4182__B2 _4181_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3556_ _3556_/A vssd1 vssd1 vccd1 vccd1 _3556_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2732__A2 _2621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4658__A _4660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3487_ _3493_/A _5639_/Q vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__and2_1
XANTENNA__3562__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput109 ksc_dat_i[0] vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__clkbuf_2
X_5226_ _5226_/A vssd1 vssd1 vccd1 vccd1 _5742_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3281__B _5533_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5157_ _5176_/A _5167_/B _5157_/C vssd1 vssd1 vccd1 vccd1 _5158_/A sky130_fd_sc_hd__or3_1
XFILLER_44_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _3932_/X _5680_/Q _4107_/Y _3934_/X vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5088_ _5081_/X _5078_/X _5087_/X _5084_/X _4026_/B vssd1 vssd1 vccd1 vccd1 _5675_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4393__A _4393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4039_ _3932_/X _5676_/Q _4038_/Y _3934_/X vssd1 vssd1 vccd1 vccd1 _4041_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3996__A1 _3996_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5639__D _5639_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3737__A _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5374__D _5374_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input174_A spi_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__A2 _4439_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3920__A1 _3794_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4568__A _5042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3903__C _3903_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4287__B _5310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A cpu_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4881__C1 _4848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2816__A _2902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4633__C1 _4632_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3411__S _3432_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5549__D _5549_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output393_A _3153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3647__A _3647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2551__A _2621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5431__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2962__A2 _2882_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3410_ _3410_/A vssd1 vssd1 vccd1 vccd1 _3410_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4164__A1 _3735_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__B_N _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4390_ _4390_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__or2_1
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2714__A2 _2621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3911__A1 _3824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3341_ _4830_/A vssd1 vssd1 vccd1 vccd1 _3357_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4478__A _4487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5581__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3382__A _3418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__C _4909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__B1 _5102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3272_ _3267_/X _3268_/X _4773_/A vssd1 vssd1 vccd1 vccd1 _3272_/X sky130_fd_sc_hd__o21a_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4219__A2 _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2726__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5102__A _5102_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5459__D _5459_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4941__A _4941_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5775_ _5800_/CLK _5775_/D vssd1 vssd1 vccd1 vccd1 _5775_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4660__B _4660_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ _5742_/Q input31/X _3246_/S vssd1 vssd1 vccd1 vccd1 _5225_/A sky130_fd_sc_hd__mux2_2
XFILLER_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4726_ _4726_/A _4731_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__and3_1
XFILLER_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4657_ _5478_/Q _4652_/X _4202_/X _4621_/A vssd1 vssd1 vccd1 vccd1 _5478_/D sky130_fd_sc_hd__a211o_1
XANTENNA__4155__A1 _5790_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput80 gpio_dat_i[15] vssd1 vssd1 vccd1 vccd1 _4048_/C sky130_fd_sc_hd__clkbuf_1
X_3608_ _3608_/A vssd1 vssd1 vccd1 vccd1 _3636_/S sky130_fd_sc_hd__buf_2
XANTENNA__4155__B2 _4154_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput91 gpio_dat_i[25] vssd1 vssd1 vccd1 vccd1 _4205_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4588_ _4588_/A vssd1 vssd1 vccd1 vccd1 _5437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3539_ _4306_/A _5596_/Q _3642_/S vssd1 vssd1 vccd1 vccd1 _4909_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4388__A _4396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3292__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5104__B1 _5097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5209_ _5209_/A vssd1 vssd1 vccd1 vccd1 _5734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4863__C1 _4843_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4554__C _4554_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5369__D _5369_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2641__A1 _2616_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5454__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4146__A1 _5474_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3914__B _5282_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4298__A _4298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4729__C _4729_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output239_A _3274_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5110__A3 _4872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3930__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4854__C1 _4840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2546__A _5767_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output406_A _3222_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4606__C1 _4598_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4464__C _4485_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2980__S _3229_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _2910_/A _2910_/B _2910_/C vssd1 vssd1 vccd1 vccd1 _2910_/Y sky130_fd_sc_hd__nor3_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4761__A _4761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3890_ _4062_/A vssd1 vssd1 vccd1 vccd1 _3890_/X sky130_fd_sc_hd__buf_4
XFILLER_91_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2841_ _2841_/A _2909_/B _2909_/C _2929_/B vssd1 vssd1 vccd1 vccd1 _2842_/C sky130_fd_sc_hd__nand4_1
XANTENNA__3377__A _3377_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5560_ _5589_/CLK _5560_/D vssd1 vssd1 vccd1 vccd1 _5560_/Q sky130_fd_sc_hd__dfxtp_1
X_2772_ _4117_/A vssd1 vssd1 vccd1 vccd1 _3331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4511_ _4511_/A vssd1 vssd1 vccd1 vccd1 _5406_/D sky130_fd_sc_hd__clkbuf_1
X_5491_ _5531_/CLK _5491_/D vssd1 vssd1 vccd1 vccd1 _5491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4442_ _4442_/A vssd1 vssd1 vccd1 vccd1 _5381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5742__D _5742_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4373_ _4373_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__or2_1
XANTENNA__3896__B1 _3886_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3324_/A vssd1 vssd1 vccd1 vccd1 _3324_/X sky130_fd_sc_hd__clkbuf_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5098__C1 _4109_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5327__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3648__A0 _4292_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4936__A _4936_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3255_ _4381_/A _5524_/Q _3444_/S vssd1 vssd1 vccd1 vccd1 _4763_/C sky130_fd_sc_hd__mux2_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__A3 _5090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3840__A _4153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4845__C1 _4840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3186_ _5724_/Q input49/X _3186_/S vssd1 vssd1 vccd1 vccd1 _5184_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2871__A1 _5694_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5477__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4671__A _4671_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4390__B _4425_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3287__A _3287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5758_ _5767_/CLK _5758_/D vssd1 vssd1 vccd1 vccd1 _5758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4709_ _4724_/A _4714_/B _4709_/C vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__or3_1
XFILLER_100_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _5690_/CLK _5689_/D vssd1 vssd1 vccd1 vccd1 _5689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5652__D _5652_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5007__A _5007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3639__A0 _4368_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4846__A _4846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3750__A _3846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input137_A ksc_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4851__A2 _3893_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2862__A1 _2809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3900__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4064__B1 _3998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4603__A2 _4589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2813__B _2831_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output189_A _4123_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4119__A1 _4114_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output356_A _3002_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5562__D _5562_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__B1 _5745_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2975__S _3233_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4756__A _4756_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3660__A _3660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4827__C1 _4823_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5095__A2 _5094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3040_ _3042_/A _5450_/Q vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__and2_1
XFILLER_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4475__B _4475_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4991_/A vssd1 vssd1 vccd1 vccd1 _5628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5252__C1 _5235_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4491__A _4491_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3942_ _3832_/X _3833_/X _3942_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _3942_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__3802__B1 _3792_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3873_ _3769_/X _3770_/X _3873_/C _4278_/D vssd1 vssd1 vccd1 vccd1 _3873_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__5737__D _5737_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5612_ _5692_/CLK _5612_/D vssd1 vssd1 vccd1 vccd1 _5612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2824_ _2806_/X _2699_/X _5375_/Q vssd1 vssd1 vccd1 vccd1 _4431_/C sky130_fd_sc_hd__a21o_2
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5543_ _5555_/CLK _5543_/D vssd1 vssd1 vccd1 vccd1 _5543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2755_ _2605_/Y _2540_/X _2794_/C _2611_/Y vssd1 vssd1 vccd1 vccd1 _2755_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5307__B1 _4240_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5474_ _5482_/CLK _5474_/D vssd1 vssd1 vccd1 vccd1 _5474_/Q sky130_fd_sc_hd__dfxtp_1
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2831_/D sky130_fd_sc_hd__clkbuf_2
X_4425_ _4425_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__or2_1
XANTENNA__5472__D _5472_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4356_ _4356_/A vssd1 vssd1 vccd1 vccd1 _5340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3307_ _3307_/A vssd1 vssd1 vccd1 vccd1 _3307_/X sky130_fd_sc_hd__clkbuf_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4666__A _4666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4287_ _4287_/A _5310_/A vssd1 vssd1 vccd1 vccd1 _4287_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3570__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__A2 _4988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _5698_/Q input67/X _3246_/S vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__mux2_2
XFILLER_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _5176_/C _5336_/Q _3192_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__mux2_8
XANTENNA__2844__A1 _5590_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2914__A _3418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4061__A3 _3994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5647__D _5647_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5382__D _5382_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3183__C _4514_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5642__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4576__A _4823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3480__A _3482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5077__A2 _4890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4295__B _4295_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4285__B1 _3866_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4824__A2 _4803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5792__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2835__A1 _2806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__A _5200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2599__B1 _5750_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3260__A1 _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5557__D _5557_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2661__A1_N _5374_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2540_ _2691_/A vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__buf_4
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4189__C _4189_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4210_ _5794_/Q _4070_/X _4200_/X _4209_/Y vssd1 vssd1 vccd1 vccd1 _5304_/A sky130_fd_sc_hd__o22ai_4
X_5190_ _5190_/A vssd1 vssd1 vccd1 vccd1 _5726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4141_ _4141_/A vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__buf_4
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4486__A _4486_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3390__A _3393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3821__C _3821_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3079__A1 _5321_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4072_ _3932_/X _5678_/Q _4071_/Y _3934_/X vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__4276__B1 _3846_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _3027_/A _5442_/Q vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__and2_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2826__A1 _2806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2734__A _2761_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4974_ _4974_/A _4997_/B _4997_/C vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__and3_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5240__A2 _5234_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3925_ _3922_/X _3723_/X _3725_/X _3924_/X vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3251__A1 _5316_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5467__D _5467_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5515__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3856_ _3851_/X _3853_/Y _5087_/A vssd1 vssd1 vccd1 vccd1 _3856_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2807_ _2806_/X _2699_/X _5381_/Q vssd1 vssd1 vccd1 vccd1 _4441_/C sky130_fd_sc_hd__a21o_2
XFILLER_101_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3787_ _3869_/A _5275_/A vssd1 vssd1 vccd1 vccd1 _3787_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3565__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5526_ _5635_/CLK _5526_/D vssd1 vssd1 vccd1 vccd1 _5526_/Q sky130_fd_sc_hd__dfxtp_1
X_2738_ _2672_/A _2699_/A _2692_/Y vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5665__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3284__B _5534_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2762__B1 _2761_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5457_ _5798_/CLK _5457_/D vssd1 vssd1 vccd1 vccd1 _5457_/Q sky130_fd_sc_hd__dfxtp_1
X_2669_ _2667_/Y _2640_/X _2668_/Y _2637_/A vssd1 vssd1 vccd1 vccd1 _4441_/B sky130_fd_sc_hd__o211ai_4
XFILLER_86_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4408_ _4600_/A vssd1 vssd1 vccd1 vccd1 _4573_/D sky130_fd_sc_hd__buf_4
XFILLER_86_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5388_ _5435_/CLK _5388_/D vssd1 vssd1 vccd1 vccd1 _5388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _5332_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4396__A _4396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2909__A _2909_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2628__B _2628_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4267__B1 _4846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__A2 _4803_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2817__A1 _2700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4019__B1 _4018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__A _5042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__A1 input68/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5377__D _5377_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__A3 _2549_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3194__B _3194_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input65_A cpu_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5298__A2 _5289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2819__A _2819_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4737__C _4741_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__B1 _3768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output221_A _3304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2808__A1 _4423_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output319_A _3585_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2808__B2 _4441_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2554__A _5382_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__B _3380_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3233__A1 input59/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__B1 _2827_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3710_/A vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4690_ _4690_/A _4707_/B _4690_/C vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__and3_1
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5688__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3641_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3385__A _3385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3572_ _3608_/A vssd1 vssd1 vccd1 vccd1 _3600_/S sky130_fd_sc_hd__buf_2
XFILLER_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2744__B1 _4437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5311_ _5801_/Q _5114_/A _5069_/X _3685_/A _5287_/A vssd1 vssd1 vccd1 vccd1 _5801_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5242_ _5266_/C _2676_/X _4848_/A vssd1 vssd1 vccd1 vccd1 _5242_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4928__B _4940_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2729__A _4617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5750__D _5750_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5173_ _5173_/A vssd1 vssd1 vccd1 vccd1 _5719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5105__A _5105_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4124_ _4196_/A vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__buf_4
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 RST_N vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XANTENNA__4944__A _5005_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4055_ _4055_/A vssd1 vssd1 vccd1 vccd1 _4055_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3006_ _3006_/A vssd1 vssd1 vccd1 vccd1 _3006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3472__A1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3279__B _5532_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4957_ _4957_/A _4965_/B _4965_/C vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__and3_1
XANTENNA__3224__A1 _5346_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3775__A2 _3756_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3908_ _4117_/A vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4888_ _3662_/Y _3678_/X _4847_/X _4271_/Y _4848_/X vssd1 vssd1 vccd1 vccd1 _5587_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__2983__A0 _5741_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3839_ _3824_/X _3825_/X _3826_/X _3838_/Y vssd1 vssd1 vccd1 vccd1 _3839_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__2911__B _2911_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3295__A _3303_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__C _2864_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__B1 _5758_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5509_ _5555_/CLK _5509_/D vssd1 vssd1 vccd1 vccd1 _5509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput360 _3011_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput371 _3033_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput382 _2990_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[7] sky130_fd_sc_hd__buf_2
Xoutput393 _3153_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__2639__A _2639_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5660__D _5660_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3234__S _3234_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5015__A _5015_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4573__B _5431_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3463__A1 _5630_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__B _3194_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3215__A1 _5414_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4191__A2 _3828_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output269_A _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3933__A _3933_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2549__A _2549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5570__D _5570_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3151__A0 _4340_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5360__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2983__S _3233_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4764__A _4764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3454__A1 _3281_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__B _4498_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _4821_/A _5545_/Q _4817_/C vssd1 vssd1 vccd1 vccd1 _4812_/A sky130_fd_sc_hd__and3_1
XANTENNA__3099__B _3105_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5791_ _5802_/CLK _5791_/D vssd1 vssd1 vccd1 vccd1 _5791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4403__B1 _4402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4742_ _4742_/A vssd1 vssd1 vccd1 vccd1 _5515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4930__C _4930_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2965__A0 _5215_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4743_/A vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__buf_4
XANTENNA__5745__D _5745_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3624_ _3630_/A _3637_/B _4965_/A vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__and3_1
XANTENNA__2717__B1 _2716_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3555_ _3558_/A _3565_/B _4920_/C vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__and3_1
XANTENNA__4182__A2 _4070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4939__A _4939_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3843__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3486_ _3486_/A vssd1 vssd1 vccd1 vccd1 _3486_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4658__B _4658_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3562__B _3565_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5225_ _5225_/A _5225_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__and3_1
XANTENNA__5480__D _5480_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5703__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5156_ _5156_/A vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4107_ _4107_/A vssd1 vssd1 vccd1 vccd1 _4107_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4674__A _4674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5087_ _5087_/A vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4038_ _4038_/A vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3996__A2 _3954_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2922__A _5660_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5655__D _5655_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3229__S _3229_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3753__A _3848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3920__A2 _3919_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input167_A spi_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5383__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5390__D _5390_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput190 _3787_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3133__A0 _4333_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4881__B1 _4191_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input28_A cpu_adr_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4584__A _4617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2816__B _2902_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4633__B1 _3878_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5565__D _5565_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output386_A _3055_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3139__S _3162_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4164__A2 _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4759__A _4759_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5726__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3372__A0 _4327_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3340_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3911__A2 _3825_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4478__B _4498_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _5099_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3271_ _4392_/B _5529_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__mux2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5056_/D vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__clkbuf_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3675__A1 _4098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4494__A _4514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4085__D1 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2986_ _2973_/X _2974_/X _4558_/C vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__o21a_1
X_5774_ _5800_/CLK _5774_/D vssd1 vssd1 vccd1 vccd1 _5774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2938__B1 _5627_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4725_ _4725_/A vssd1 vssd1 vccd1 vccd1 _5508_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5475__D _5475_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4656_ _3756_/X _4667_/C _4186_/Y _4185_/X _4630_/X vssd1 vssd1 vccd1 vccd1 _5477_/D
+ sky130_fd_sc_hd__o221a_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__clkbuf_1
Xinput70 cpu_sel_i[3] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_2
Xinput81 gpio_dat_i[16] vssd1 vssd1 vccd1 vccd1 _4063_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__4155__A2 _4070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4587_ _4592_/A _5437_/Q _4604_/C _4596_/D vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__and4_1
XANTENNA__4669__A _4746_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput92 gpio_dat_i[26] vssd1 vssd1 vccd1 vccd1 _4217_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3538_ _3608_/A vssd1 vssd1 vccd1 vccd1 _3642_/S sky130_fd_sc_hd__buf_4
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__B _4388_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3292__B _5538_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5104__A1 _5096_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3469_ _3530_/A vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__A0 _5154_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5208_ _5208_/A _5225_/B _5208_/C vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__and3_1
XFILLER_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4863__B1 _4856_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5139_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5705_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2917__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__B _2761_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2641__A2 _2617_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3748__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2652__A _2652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5385__D _5385_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5749__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4146__A2 _4074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4579__A _4592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3483__A _3483_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3657__A1 _3711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4854__B1 _3944_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3930__B _3930_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3422__S _3435_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5203__A _5203_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4606__B1 _3062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output301_A _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4761__B _4778_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2840_ _2839_/Y _2762_/Y _4411_/C vssd1 vssd1 vccd1 vccd1 _2929_/B sky130_fd_sc_hd__a21oi_2
X_2771_ _2771_/A vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__buf_2
XANTENNA__3593__A0 _4340_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4510_ _4514_/A _4524_/B _4510_/C vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__or3_1
XFILLER_34_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5490_ _5538_/CLK _5490_/D vssd1 vssd1 vccd1 vccd1 _5490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4441_ _4441_/A _4441_/B _4441_/C vssd1 vssd1 vccd1 vccd1 _4442_/A sky130_fd_sc_hd__and3_1
XANTENNA__4489__A _4489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__A _3393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4372_ _4372_/A vssd1 vssd1 vccd1 vccd1 _5347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3896__A1 _5775_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3896__B2 _3895_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3323_ _3325_/A _5552_/Q vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__and2_1
XFILLER_99_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__B1 _5097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3403_/A vssd1 vssd1 vccd1 vccd1 _3444_/S sky130_fd_sc_hd__buf_2
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3648__A1 _5591_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4936__B _4940_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__B1 _3838_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3185_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2608__B1_N _5747_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2871__A2 _4968_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4952__A _4952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4671__B _4681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3568__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _5738_/Q input27/X _3246_/S vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__mux2_2
X_5757_ _5765_/CLK _5757_/D vssd1 vssd1 vccd1 vccd1 _5757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4708_ _4708_/A vssd1 vssd1 vccd1 vccd1 _5501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5688_ _5690_/CLK _5688_/D vssd1 vssd1 vccd1 vccd1 _5688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4399__A _5195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4639_ _4652_/A vssd1 vssd1 vccd1 vccd1 _4639_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5007__B _5130_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3639__A1 _5624_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2647__A _2647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3242__S _3250_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5023__A _5097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5421__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__D1 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2862__A2 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4064__A1 _3922_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4129__B1_N _5473_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5571__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2813__C _2813_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input95_A gpio_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4119__A2 _4115_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output251_A _3394_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output349_A _3653_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3941__A _5566_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2550__A1 _2707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4756__B _4756_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4827__B1 _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5095__A3 _5087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2557__A _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4475__C _4485_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4772__A _4772_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4990_ _4990_/A _4990_/B _4990_/C vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__or3_1
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5252__B1 _2687_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4491__B _4500_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3941_ _5566_/Q vssd1 vssd1 vccd1 vccd1 _3941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3802__A1 _5771_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3388__A _3388_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3802__B2 _3801_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3872_ _5562_/Q vssd1 vssd1 vccd1 vccd1 _3872_/Y sky130_fd_sc_hd__inv_2
X_5611_ _5692_/CLK _5611_/D vssd1 vssd1 vccd1 vccd1 _5611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2823_ _2809_/X _2750_/X _5380_/Q vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_34_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5542_ _5555_/CLK _5542_/D vssd1 vssd1 vccd1 vccd1 _5542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2754_ _2569_/X _2544_/B _2549_/X _2753_/X vssd1 vssd1 vccd1 vccd1 _2794_/C sky130_fd_sc_hd__a31oi_2
XFILLER_34_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5307__A1 _5797_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5307__B2 _4247_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5473_ _5737_/CLK _5473_/D vssd1 vssd1 vccd1 vccd1 _5473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5753__D _5753_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2685_ _2761_/C vssd1 vssd1 vccd1 vccd1 _2813_/C sky130_fd_sc_hd__buf_2
X_4424_ _4424_/A vssd1 vssd1 vccd1 vccd1 _5371_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4012__A _5570_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4355_ _4355_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__or2_1
XANTENNA__4947__A _4947_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4225__A2_N _5688_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3851__A _4254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3306_ _3314_/A _5544_/Q vssd1 vssd1 vccd1 vccd1 _3307_/A sky130_fd_sc_hd__and2_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5444__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _5289_/A _5800_/Q _4282_/Y _4285_/Y vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__o22ai_4
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4279__D1 _3836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3570__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3237_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3237_/X sky130_fd_sc_hd__clkbuf_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3168_ _5721_/Q input45/X _3168_/S vssd1 vssd1 vccd1 vccd1 _5176_/C sky130_fd_sc_hd__mux2_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2844__A2 _4115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5594__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4682__A _4682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3099_ _3123_/A _3105_/B _4478_/C vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__and3_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5243__B1 _5242_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3298__A _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3557__A0 _4318_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5663__D _5663_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5018__A _5018_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4857__A _5087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3761__A _4692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3480__B _5636_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5077__A3 _5070_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4285__A1 _3707_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4295__C _4295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A cpu_adr_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2835__A2 _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4592__A _4592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2599__A1 _2616_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__B1 _3795_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5200__B _5215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3260__A2 _2899_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3001__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5317__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output299_A _3519_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3936__A _4109_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5573__D _5573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5467__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4189__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4767__A _4771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3671__A _3699_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4140_ _4140_/A vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3390__B _3397_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _4071_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4276__A1 _5692_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4276__B2 _5112_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3022_ _3022_/A vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2826__A2 _5266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4028__A1 _4027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4973_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4997_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__5748__D _5748_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2734__B _2761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4007__A _4153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3924_ _3727_/X _3729_/X _3924_/C _4063_/D vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__and4bb_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3855_ _4846_/A vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__buf_6
XANTENNA__3539__A0 _4306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3846__A _3846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2750__A _2750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2806_ _2806_/A vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__clkbuf_4
X_3786_ _3747_/X _5770_/Q _3776_/Y _3785_/Y vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__3565__B _3565_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5525_ _5531_/CLK _5525_/D vssd1 vssd1 vccd1 vccd1 _5525_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _5373_/Q _2565_/A _4427_/B vssd1 vssd1 vccd1 vccd1 _2779_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__5483__D _5483_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3057__S _3108_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2762__A1 _5746_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2668_ _2616_/X _2549_/A _5766_/Q vssd1 vssd1 vccd1 vccd1 _2668_/Y sky130_fd_sc_hd__o21ai_2
X_5456_ _5482_/CLK _5456_/D vssd1 vssd1 vccd1 vccd1 _5456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__buf_2
XANTENNA__4677__A _4677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3581__A _3594_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5387_ _5435_/CLK _5387_/D vssd1 vssd1 vccd1 vccd1 _5387_/Q sky130_fd_sc_hd__dfxtp_1
X_2599_ _2616_/A _2549_/A _5750_/Q vssd1 vssd1 vccd1 vccd1 _2600_/C sky130_fd_sc_hd__o21ai_1
XFILLER_87_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4338_ _4338_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__or2_1
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2909__B _2909_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4396__B _4396_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input2_A cpu_adr_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4269_ _3860_/X _3861_/X _4269_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__and4bb_1
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4267__A1 _4265_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2628__C _2628_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2817__A2 _5266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2925__A _2925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4019__A1 _5466_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5658__D _5658_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__B1 _4617_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3756__A _3857_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2660__A _2660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5393__D _5393_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3194__C _4520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input58_A cpu_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4587__A _4592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3491__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2819__B _2848_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__A1 _3763_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2808__A2 _4423_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output214_A _3289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5211__A _5211_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5568__D _5568_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__C _4705_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__A1 _5374_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3666__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3640_ _3646_/A _4988_/B _4980_/C vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__and3_1
XFILLER_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4194__B1 _4193_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3571_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3571_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2744__A1 _5379_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5310_ _5310_/A _5310_/B vssd1 vssd1 vccd1 vccd1 _5800_/D sky130_fd_sc_hd__nand2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4497__A _4497_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5241_ _2592_/Y _5227_/X _2595_/Y _5228_/X _4429_/X vssd1 vssd1 vccd1 vccd1 _5749_/D
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__3605__S _3633_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4928__C _4940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5172_ _5176_/A _5191_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__or3_1
XFILLER_9_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4123_ _4123_/A _5297_/A vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5105__B _5111_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput2 cpu_adr_i[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
X_4054_ _4123_/A _5293_/A vssd1 vssd1 vccd1 vccd1 _4054_/Y sky130_fd_sc_hd__nor2_8
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3005_ _3005_/A _5434_/Q vssd1 vssd1 vccd1 vccd1 _3006_/A sky130_fd_sc_hd__and2_1
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3472__A2 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5121__A _5121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2680__B1 _5752_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5478__D _5478_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4960__A _4960_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4956_ _4956_/A vssd1 vssd1 vccd1 vccd1 _5614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5632__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3907_ _3832_/X _3833_/X _3907_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__and4bb_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4887_ _4875_/X _4876_/X _4259_/Y _4877_/X vssd1 vssd1 vccd1 vccd1 _5586_/D sky130_fd_sc_hd__a211o_1
XANTENNA__2983__A1 input30/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3838_ _3827_/Y _3828_/X _3837_/Y vssd1 vssd1 vccd1 vccd1 _3838_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2911__C _2925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3295__B _5539_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__A_N _5768_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3769_ _3999_/A vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5782__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2735__A1 _2607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5508_ _5635_/CLK _5508_/D vssd1 vssd1 vccd1 vccd1 _5508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput350 _3655_/X vssd1 vssd1 vccd1 vccd1 ksc_sel_o[3] sky130_fd_sc_hd__buf_2
X_5439_ _5446_/CLK _5439_/D vssd1 vssd1 vccd1 vccd1 _5439_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput361 _3013_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_82_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput372 _3035_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput383 _2993_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[8] sky130_fd_sc_hd__buf_2
XANTENNA__4200__A _4252_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput394 _3160_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3250__S _3250_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5031__A _5043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4573__C _4665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input112_A ksc_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5388__D _5388_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__C _4517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4056__A2_N _5677_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3486__A _3486_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3425__S _3432_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5206__A _5206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4110__A _4110_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3151__A1 _5403_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5505__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output331_A _3625_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2565__A _2565_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4483__C _4483_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3454__A2 _2899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5655__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2662__B1 _2661_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _5544_/Q _4803_/X _4798_/X _4804_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5544_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4780__A _4803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3099__C _4478_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4403__A1 _2752_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5790_ _5798_/CLK _5790_/D vssd1 vssd1 vccd1 vccd1 _5790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4741_ _4741_/A _4756_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__and3_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2965__A1 _5352_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_19_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5694_/CLK sky130_fd_sc_hd__clkbuf_16
X_4672_ _4672_/A vssd1 vssd1 vccd1 vccd1 _5487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4167__B1 _4159_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3623_ _4357_/B _5619_/Q _3636_/S vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2717__A1 _2715_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ _4316_/A _5600_/Q _3642_/S vssd1 vssd1 vccd1 vccd1 _4920_/C sky130_fd_sc_hd__mux2_1
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3843__B _5277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5116__C1 _4883_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3485_ _3493_/A _5638_/Q vssd1 vssd1 vccd1 vccd1 _3486_/A sky130_fd_sc_hd__and2_1
XANTENNA__5761__D _5761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3562__C _4926_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5224_ _5224_/A vssd1 vssd1 vccd1 vccd1 _5741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4955__A _4963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5155_ _5155_/A vssd1 vssd1 vccd1 vccd1 _5712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _4123_/A _4106_/B vssd1 vssd1 vccd1 vccd1 _4106_/Y sky130_fd_sc_hd__nor2_8
X_5086_ _5674_/Q _4988_/A _3750_/X _5086_/B2 _5064_/A vssd1 vssd1 vccd1 vccd1 _5674_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4674__B _4688_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _4196_/A vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__buf_8
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3070__S _3108_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2653__B1 _5762_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3996__A3 _3994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__A _4690_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _5608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4158__B1 _4157_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3972__B_N _3818_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5107__C1 _4214_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5528__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5671__D _5671_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5026__A _5033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput180 _3966_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput191 _4137_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__3133__A1 _5400_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4865__A _5235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4881__A1 _3662_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5678__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2892__B1 _3073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4633__A1 _5458_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2816__C _2816_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2644__B1 _2544_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3841__C1 _3840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output281_A _2915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output379_A _2978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3372__A1 _5501_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_3_0_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_1_CLK/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5581__D _5581_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3155__S _3168_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4478__C _4478_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _3267_/X _3268_/X _4771_/C vssd1 vssd1 vccd1 vccd1 _3270_/X sky130_fd_sc_hd__o21a_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A2 _5094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4775__A _4917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3675__A2 _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5446_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2883__B1 _5266_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4494__B _4498_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4085__C1 _4084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5756__D _5756_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5773_ _5802_/CLK _5773_/D vssd1 vssd1 vccd1 vccd1 _5773_/Q sky130_fd_sc_hd__dfxtp_1
X_2985_ _4394_/A _5426_/Q _3252_/S vssd1 vssd1 vccd1 vccd1 _4558_/C sky130_fd_sc_hd__mux2_1
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2938__A1 _2929_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4724_ _4724_/A _4739_/B _4724_/C vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__or3_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4655_ _5476_/Q _4652_/X _4174_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _5476_/D sky130_fd_sc_hd__a211o_1
XFILLER_11_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3606_ _3613_/A _3620_/B _4955_/C vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__and3_1
Xinput60 cpu_dat_i[3] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput71 cpu_stb_i vssd1 vssd1 vccd1 vccd1 _2581_/A sky130_fd_sc_hd__buf_6
X_4586_ _5042_/A vssd1 vssd1 vccd1 vccd1 _4604_/C sky130_fd_sc_hd__clkbuf_2
Xinput82 gpio_dat_i[17] vssd1 vssd1 vccd1 vccd1 _4084_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput93 gpio_dat_i[27] vssd1 vssd1 vccd1 vccd1 _4231_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3537_ _3537_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5491__D _5491_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3065__S _5234_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5104__A2 _5089_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3468_ _2924_/X _2927_/X _4997_/A vssd1 vssd1 vccd1 vccd1 _3468_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__A1 _5327_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4685__A _4711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3399_ _3418_/A vssd1 vssd1 vccd1 vccd1 _3416_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4863__A1 _4002_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4863__B2 _4857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5138_ _5152_/A _5143_/B _5138_/C vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__or3_1
XANTENNA__2917__B _2917_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__buf_4
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__C _2647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5666__D _5666_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5350__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3764__A _3980_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4579__B _5433_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2562__C1 _2561_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A cpu_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4595__A _4595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3657__A2 _2854_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4854__A1 _4836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4606__A1 _5446_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4067__C1 _4007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4606__B2 _4590_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3004__A _3004_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4761__C _4765_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5576__D _5576_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _3736_/A vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__inv_2
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3593__A1 _5611_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2989__S _3240_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3674__A _3674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4440_ _4440_/A vssd1 vssd1 vccd1 vccd1 _5380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3393__B _3397_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4371_ _4396_/A _4371_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__and2_1
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3896__A2 _3690_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3322_ _3322_/A vssd1 vssd1 vccd1 vccd1 _3322_/X sky130_fd_sc_hd__clkbuf_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4001__C _4001_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A1 _5096_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _2994_/A _2882_/A _4456_/C vssd1 vssd1 vccd1 vccd1 _3253_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4936__C _4940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__A1 _4836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3184_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3184_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2856__B1 _4617_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3849__A _3849_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2753__A _5556_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4671__C _4690_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5486__D _5486_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5373__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5756_ _5767_/CLK _5756_/D vssd1 vssd1 vccd1 vccd1 _5756_/Q sky130_fd_sc_hd__dfxtp_1
X_2968_ _3179_/A vssd1 vssd1 vccd1 vccd1 _3246_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4707_ _4707_/A _4707_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__and3_1
XANTENNA__4173__B_N _4076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5687_ _5690_/CLK _5687_/D vssd1 vssd1 vccd1 vccd1 _5687_/Q sky130_fd_sc_hd__dfxtp_1
X_2899_ _2899_/A vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3584__A _3594_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2792__C1 _2540_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4638_ _4638_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _5463_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _4569_/A _5429_/Q _4665_/D _4573_/D vssd1 vssd1 vccd1 vccd1 _4570_/A sky130_fd_sc_hd__and4_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5007__C _5021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5304__A _5304_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__B1 _5360_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4049__C1 _4048_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5246__D1 _5236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4064__A2 _3958_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5716__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3759__A _5558_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2663__A _2761_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3272__B1 _4773_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5396__D _5396_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2813__D _2831_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4221__C1 _3840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input88_A gpio_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__A _3494_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__A2 _2549_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output244_A _3336_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4827__A1 _5554_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4756__C _4765_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5214__A _5214_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4827__B2 _4804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2838__B1 _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2557__B _2583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output411_A _3074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5237__D1 _5236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5396__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5252__A1 _5758_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__A _4665_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2573__A _2573_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3940_ _4147_/A vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4491__C _4512_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3802__A2 _3690_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _5666_/Q _5002_/A _3846_/X _5073_/B2 vssd1 vssd1 vccd1 vccd1 _3871_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5610_ _5692_/CLK _5610_/D vssd1 vssd1 vccd1 vccd1 _5610_/Q sky130_fd_sc_hd__dfxtp_1
X_2822_ _2817_/X _2642_/Y _2821_/Y vssd1 vssd1 vccd1 vccd1 _2902_/B sky130_fd_sc_hd__a21oi_4
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5541_ _5555_/CLK _5541_/D vssd1 vssd1 vccd1 vccd1 _5541_/Q sky130_fd_sc_hd__dfxtp_1
X_2753_ _5556_/Q _5696_/Q vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__or2_1
XFILLER_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3835__C _3835_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5307__A2 _5268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5472_ _5798_/CLK _5472_/D vssd1 vssd1 vccd1 vccd1 _5472_/Q sky130_fd_sc_hd__dfxtp_1
X_2684_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2831_/B sky130_fd_sc_hd__clkbuf_2
X_4423_ _4431_/A _4423_/B _4423_/C vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__and3_1
XFILLER_82_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4354_ _4354_/A vssd1 vssd1 vccd1 vccd1 _5339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3851__B _4265_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3305_ _3316_/A vssd1 vssd1 vccd1 vccd1 _3314_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2748__A _2782_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4285_ _3707_/X _4284_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _4285_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4279__C1 _4278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5124__A _5128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3570__C _4930_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3236_/A _4542_/B _4538_/C vssd1 vssd1 vccd1 vccd1 _3237_/A sky130_fd_sc_hd__and3_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5739__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4963__A _4963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3167_ _3196_/A vssd1 vssd1 vccd1 vccd1 _3194_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3098_ _4320_/A _5394_/Q _3146_/S vssd1 vssd1 vccd1 vccd1 _4478_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5243__A1 _2600_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3579__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3557__A1 _5601_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5739_ _5741_/CLK _5739_/D vssd1 vssd1 vccd1 vccd1 _5739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2765__C1 _2691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5034__A _5034_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input142_A ksc_rty_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4285__A2 _4284_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4295__D _4295_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4873__A _5087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4592__B _5439_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3489__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3245__B1 _4451_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2599__A2 _2549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__A1 _3796_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__C _5200_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_1_1_CLK_A clkbuf_opt_1_1_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3001__B _5432_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3936__B _3936_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output194_A _4183_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3428__S _3435_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5209__A _5209_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output361_A _3013_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4767__B _4776_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4160__B1_N _5475_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3671__B _3698_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2568__A _5382_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3390__C _4719_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4070_/A vssd1 vssd1 vccd1 vccd1 _4070_/X sky130_fd_sc_hd__buf_4
XFILLER_42_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4276__A2 _5002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3021_ _3027_/A _5441_/Q vssd1 vssd1 vccd1 vccd1 _3022_/A sky130_fd_sc_hd__and2_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4783__A _4823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4028__A2 _3919_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3399__A _3418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4972_ _5183_/A vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_52_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4433__C1 _2783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2734__C _2734_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3923_ _4099_/A vssd1 vssd1 vccd1 vccd1 _4063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3854_ _2845_/X _4128_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__o21a_4
XANTENNA__3539__A1 _5596_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2805_ _2569_/X _2559_/X _5371_/Q vssd1 vssd1 vccd1 vccd1 _4423_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5764__D _5764_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3785_ _5089_/A _3783_/Y _5289_/A vssd1 vssd1 vccd1 vccd1 _3785_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3338__S _3441_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5119__A _5212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3565__C _4928_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5524_ _5635_/CLK _5524_/D vssd1 vssd1 vccd1 vccd1 _5524_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4023__A _4023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2736_ _2736_/A _2736_/B _2736_/C vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__nand3_2
XANTENNA__5411__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2762__A2 _2785_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5455_ _5741_/CLK _5455_/D vssd1 vssd1 vccd1 vccd1 _5455_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4958__A _4958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2667_ _2667_/A vssd1 vssd1 vccd1 vccd1 _2667_/Y sky130_fd_sc_hd__clkinv_2
X_4406_ _4406_/A vssd1 vssd1 vccd1 vccd1 _5362_/D sky130_fd_sc_hd__clkbuf_1
X_5386_ _5435_/CLK _5386_/D vssd1 vssd1 vccd1 vccd1 _5386_/Q sky130_fd_sc_hd__dfxtp_1
X_2598_ _2647_/A _2686_/A input8/X _2684_/A vssd1 vssd1 vccd1 vccd1 _2600_/B sky130_fd_sc_hd__nand4_2
XANTENNA__3581__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4337_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5561__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2909__C _2909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _5587_/Q vssd1 vssd1 vccd1 vccd1 _4268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4267__A2 _4266_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4693__A _4776_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3475__A0 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3219_ _5198_/A _5345_/Q _3219_/S vssd1 vssd1 vccd1 vccd1 _4366_/B sky130_fd_sc_hd__mux2_8
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2925__B _2925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4019__A2 _4444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3778__A1 _2561_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2941__A _3622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5674__D _5674_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3248__S _3248_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5029__A _5058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4587__B _5437_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3491__B _5641_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2819__C _2848_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__A2 _3766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4663__C1 _4621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3218__A0 _5730_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output207_A _3897_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3012__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__A2 _4429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5434__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5584__D _5584_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3158__S _3204_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4194__A1 _5793_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3570_ _3577_/A _3584_/B _4930_/C vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__and3_1
XFILLER_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4239__A2_N _5689_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2744__A2 _2613_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4778__A _4778_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5584__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3682__A _3682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5240_ _5748_/Q _5234_/X _2585_/Y _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5748_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5171_ _5223_/B vssd1 vssd1 vccd1 vccd1 _5191_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4122_ _5788_/Q _4070_/X _4109_/X _4121_/Y vssd1 vssd1 vccd1 vccd1 _5297_/A sky130_fd_sc_hd__o22ai_4
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3457__A0 _4381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4053_ _5784_/Q _3804_/X _4041_/X _4052_/Y vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__o22ai_4
Xinput3 cpu_adr_i[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3004_ _3004_/A vssd1 vssd1 vccd1 vccd1 _3004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5759__D _5759_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3209__A0 _4362_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2680__A1 _2593_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4018__A _4283_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4955_ _4963_/A _4963_/B _4955_/C vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__or3_1
XANTENNA__3857__A _3857_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2761__A _2761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3906_ _4692_/A vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ _4244_/X _4245_/X _4872_/X _4873_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _5585_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5494__D _5494_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3837_ _3829_/X _3830_/X _3831_/X _3835_/X _3836_/X vssd1 vssd1 vccd1 vccd1 _3837_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2911__D _2925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3768_ _3768_/A vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5507_ _5635_/CLK _5507_/D vssd1 vssd1 vccd1 vccd1 _5507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2735__A2 _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4688__A _4699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2719_ _2719_/A vssd1 vssd1 vccd1 vccd1 _2831_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__3592__A _3592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3699_ _3697_/X _3699_/B _5034_/A vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__nand3b_4
X_5438_ _5446_/CLK _5438_/D vssd1 vssd1 vccd1 vccd1 _5438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput340 _3548_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput351 _5806_/X vssd1 vssd1 vccd1 vccd1 ksc_stb_o sky130_fd_sc_hd__buf_2
XFILLER_86_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput362 _3015_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput373 _3037_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[28] sky130_fd_sc_hd__buf_2
XFILLER_82_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput384 _2995_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5369_ _5695_/CLK _5369_/D vssd1 vssd1 vccd1 vccd1 _5369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4200__B _4200_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput395 _3166_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[18] sky130_fd_sc_hd__buf_2
XANTENNA__4893__C1 _4630_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3448__B1 _4671_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5669__D _5669_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5031__B _5645_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4573__D _4573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5457__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input105_A gpio_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__A _3979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4257__B_N _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input70_A cpu_sel_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4598__A _4823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3007__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4884__C1 _4883_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output324_A _3602_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3441__S _3441_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5222__A _5222_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5579__D _5579_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2662__A1 _2657_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4403__A2 _2552_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4740_ _4740_/A vssd1 vssd1 vccd1 vccd1 _5514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2581__A _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4671_ _4671_/A _4681_/B _4690_/C vssd1 vssd1 vccd1 vccd1 _4672_/A sky130_fd_sc_hd__and3_1
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4167__A1 _5791_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3622_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3637_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4167__B2 _4166_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2717__A2 _2640_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3553_ _3553_/A vssd1 vssd1 vccd1 vccd1 _3553_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3616__S _3636_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5116__B1 _4667_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4301__A _4301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3484_ _3530_/A vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5223_ _5223_/A _5223_/B _5223_/C vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__or3_1
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5154_ _5154_/A _5154_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5155_/A sky130_fd_sc_hd__and3_1
XANTENNA__4955__B _4963_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _5787_/Q _4091_/X _4094_/X _4104_/Y vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__o22ai_4
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5081_/X _5078_/X _5066_/X _5084_/X _3993_/B vssd1 vssd1 vccd1 vccd1 _5673_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4627__C1 _4660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4674__C _4674_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5132__A _5156_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A _4036_/B vssd1 vssd1 vccd1 vccd1 _4036_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5489__D _5489_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4971__A _4971_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2653__A1 _2607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__B _4707_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5052__C1 _5045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4938_ _4938_/A _4938_/B _4938_/C vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__or3_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4869_ _4859_/X _4860_/X _4086_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5574_/D sky130_fd_sc_hd__a211o_1
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4158__B2 _3808_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5107__B1 _5102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4211__A _4263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput181 _3987_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput192 _4156_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[21] sky130_fd_sc_hd__buf_2
XANTENNA__4866__C1 _4865_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4881__A2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2892__A1 _2876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3261__S _3444_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5042__A _5042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5399__D _5399_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2816__D _2816_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4633__A2 _4623_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2644__A1 _5261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3841__B1 _3839_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3497__A _3497_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3797__B_N _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output274_A _3366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5217__A _5217_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A3 _5066_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5622__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2576__A _5261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2883__A1 _2544_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4494__C _4494_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4084__A_N _4082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4085__B1 _3979_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4791__A _4791_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5772__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5772_ _5800_/CLK _5772_/D vssd1 vssd1 vccd1 vccd1 _5772_/Q sky130_fd_sc_hd__dfxtp_1
X_2984_ _5223_/C _5356_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__mux2_8
XANTENNA__3200__A _3210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4723_ _4723_/A vssd1 vssd1 vccd1 vccd1 _5507_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2938__A2 _2937_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4654_ _4660_/A _4654_/B vssd1 vssd1 vccd1 vccd1 _5475_/D sky130_fd_sc_hd__nor2_1
X_3605_ _4346_/A _5614_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _4955_/C sky130_fd_sc_hd__mux2_1
XFILLER_11_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 cpu_dat_i[23] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 cpu_dat_i[4] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
X_4585_ _5436_/Q _4563_/X _4584_/X _4564_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _5436_/D
+ sky130_fd_sc_hd__a221o_1
Xinput72 cpu_we_i vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_2
XANTENNA__5772__D _5772_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3899__B1 _3898_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput83 gpio_dat_i[18] vssd1 vssd1 vccd1 vccd1 _4100_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5127__A _5127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput94 gpio_dat_i[28] vssd1 vssd1 vccd1 vccd1 _4243_/C sky130_fd_sc_hd__clkbuf_1
X_3536_ _3540_/A _3547_/B _4907_/A vssd1 vssd1 vccd1 vccd1 _3537_/A sky130_fd_sc_hd__and3_1
XANTENNA__2571__B1 _2570_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3467_ _4388_/B _5631_/Q _3652_/S vssd1 vssd1 vccd1 vccd1 _4997_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4966__A _4966_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3870__A _4287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5104__A3 _5090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5206_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5733_/D sky130_fd_sc_hd__clkbuf_1
X_3398_ _3398_/A vssd1 vssd1 vccd1 vccd1 _3398_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4863__A2 _4004_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5137_ _5137_/A vssd1 vssd1 vccd1 vccd1 _5704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2917__C _2917_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__buf_2
XFILLER_96_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2636__D _2761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4019_ _5466_/Q _4444_/A _4018_/X vssd1 vssd1 vccd1 vccd1 _4019_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5682__D _5682_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5037__A _5037_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4579__C _4665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input172_A spi_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5645__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2562__B1 _2560_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4876__A _5089_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3780__A _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A cpu_adr_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4854__A2 _4837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5795__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4067__B1 _4066_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4606__A2 _4589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5016__C1 _4823_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3020__A _3020_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output391_A _3142_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3674__B _3682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5592__D _5592_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__C _4722_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4370_ _4378_/A vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2553__B1 _2552_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3321_ _3325_/A _5551_/Q vssd1 vssd1 vccd1 vccd1 _3322_/A sky130_fd_sc_hd__and2_1
XANTENNA__4786__A _4828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3690__A _4091_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4001__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A2 _5089_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3252_ _4301_/A _5386_/Q _3252_/S vssd1 vssd1 vccd1 vccd1 _4456_/C sky130_fd_sc_hd__mux2_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__A2 _4837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3183_/A _3194_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _3184_/A sky130_fd_sc_hd__and3_1
XANTENNA__2856__A1 _2561_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2608__A1 _2607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5767__D _5767_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2753__B _5696_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5518__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4026__A _4127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5755_ _5800_/CLK _5755_/D vssd1 vssd1 vccd1 vccd1 _5755_/Q sky130_fd_sc_hd__dfxtp_1
X_2967_ _2876_/X _2882_/X _4550_/C vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__o21a_1
X_4706_ _4706_/A vssd1 vssd1 vccd1 vccd1 _5500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5668__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5686_ _5690_/CLK _5686_/D vssd1 vssd1 vccd1 vccd1 _5686_/Q sky130_fd_sc_hd__dfxtp_1
X_2898_ _4295_/C vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__buf_2
XANTENNA__3584__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2792__B1 _2791_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3675__B1_N _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4637_ _5462_/Q _4623_/X _3938_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _5462_/D sky130_fd_sc_hd__a211o_1
XFILLER_85_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4568_ _5042_/A vssd1 vssd1 vccd1 vccd1 _4665_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3519_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3741__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4696__A _4778_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4499_ _4499_/A vssd1 vssd1 vccd1 vccd1 _5402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5304__B _5308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__A1 _2809_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3105__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4049__B1 _3979_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5246__C1 _5235_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2944__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3272__A1 _3267_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2663__B _2761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5677__D _5677_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_0_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_1_CLK/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4221__B1 _4220_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2783__B1 _5761_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3835__B_N _3833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4827__A2 _4803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output237_A _3270_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2838__A1 _2835_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3015__A _3015_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5237__C1 _5235_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2854__A _3709_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output404_A _3211_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5252__A2 _5234_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__B _3669_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5587__D _5587_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3870_ _4287_/A vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__buf_8
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4072__A1_N _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2821_ _2818_/Y _2540_/X _2820_/Y vssd1 vssd1 vccd1 vccd1 _2821_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_73_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3685__A _3685_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5540_ _5555_/CLK _5540_/D vssd1 vssd1 vccd1 vccd1 _5540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2752_ _2675_/A _2750_/X _2751_/Y vssd1 vssd1 vccd1 vccd1 _2752_/Y sky130_fd_sc_hd__o21ai_2
X_5471_ _5737_/CLK _5471_/D vssd1 vssd1 vccd1 vccd1 _5471_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3835__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2683_ _2785_/A vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4422_ _4422_/A vssd1 vssd1 vccd1 vccd1 _5370_/D sky130_fd_sc_hd__clkbuf_1
X_5803__424 vssd1 vssd1 vccd1 vccd1 _5803__424/HI cpu_err_o sky130_fd_sc_hd__conb_1
XFILLER_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _4366_/A _4353_/B vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__and2_1
XFILLER_82_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__clkbuf_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3851__C _4283_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _5484_/Q _4444_/A _4283_/X vssd1 vssd1 vccd1 vccd1 _4284_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_87_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2748__B _2748_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4279__B1 _3768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5124__B _5143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _4373_/A _5418_/Q _3235_/S vssd1 vssd1 vccd1 vccd1 _4538_/C sky130_fd_sc_hd__mux2_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3166_ _3166_/A vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4963__B _4963_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5340__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3097_ _3163_/A vssd1 vssd1 vccd1 vccd1 _3146_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__5140__A _5264_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5243__A2 _2600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5497__D _5497_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5490__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5807_ _5807_/A vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4203__B1 _4202_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3999_ _3999_/A vssd1 vssd1 vccd1 vccd1 _3999_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3595__A _3595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5738_ _5765_/CLK _5738_/D vssd1 vssd1 vccd1 vccd1 _5738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2765__B1 _2764_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5697_/CLK _5669_/D vssd1 vssd1 vccd1 vccd1 _5669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__B _2695_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A ksc_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2674__A _2748_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__A _5056_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4592__C _4604_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3489__B _5640_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3245__A1 _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__A2 _4528_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3936__C _4240_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2756__B1 _2755_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output187_A _4090_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output354_A _2998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3444__S _3444_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3181__A0 _5181_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4767__C _4767_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5225__A _5225_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__B_N _3861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5363__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _3020_/A vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2584__A _2686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _4971_/A vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__buf_12
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4433__B1 _5238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2734__D _2761_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3922_ _4098_/A vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3853_ _2728_/A _4590_/A _5457_/Q vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3619__S _3633_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2804_ _2650_/A _2650_/B _4425_/A vssd1 vssd1 vccd1 vccd1 _2902_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__4304__A _4322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3784_ _4070_/A vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__buf_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5523_ _5538_/CLK _5523_/D vssd1 vssd1 vccd1 vccd1 _5523_/Q sky130_fd_sc_hd__dfxtp_1
X_2735_ _2607_/X _2708_/A _5758_/Q vssd1 vssd1 vccd1 vccd1 _2736_/C sky130_fd_sc_hd__o21ai_1
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5454_ _5482_/CLK _5454_/D vssd1 vssd1 vccd1 vccd1 _5454_/Q sky130_fd_sc_hd__dfxtp_1
X_2666_ _5371_/Q _2611_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _2779_/A sky130_fd_sc_hd__o21ai_4
XFILLER_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4405_ _4405_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__or2_1
XFILLER_47_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5385_ _5435_/CLK _5385_/D vssd1 vssd1 vccd1 vccd1 _5385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5706__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2759__A _2916_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5780__D _5780_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2597_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2637_/A sky130_fd_sc_hd__buf_4
XANTENNA__5135__A _5183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3581__C _4936_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4336_ _4336_/A vssd1 vssd1 vccd1 vccd1 _5331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2909__D _2929_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4974__A _4974_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4267_ _4265_/X _4266_/Y _4846_/A vssd1 vssd1 vccd1 vccd1 _4267_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4121__C1 _3946_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3218_ _5730_/Q input55/X _3228_/S vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3475__A1 _5634_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4198_ _4139_/X _5686_/Q _4197_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3149_ _5718_/Q input42/X _3186_/S vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__mux2_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2925__C _2925_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3778__A2 _3157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2986__B1 _4558_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4214__A _4240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2738__B1 _2692_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5386__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5690__D _5690_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4587__C _4604_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5045__A _5097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2819__D _2848_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4663__B1 _4283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3218__A1 input55/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3012__B _5437_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2977__A0 _4390_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4124__A _4196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4194__A2 _3690_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5729__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4778__B _4778_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2579__A _5261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5170_ _5170_/A vssd1 vssd1 vccd1 vccd1 _5718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4121_ _4042_/X _4113_/Y _4120_/Y _3946_/X vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__4794__A _4794_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4103__C1 _4005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4052_ _4042_/X _4045_/Y _4051_/Y _3946_/X vssd1 vssd1 vccd1 vccd1 _4052_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3457__A1 _5628_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 cpu_adr_i[11] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3005_/A _5433_/Q vssd1 vssd1 vccd1 vccd1 _3004_/A sky130_fd_sc_hd__and2_1
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3209__A1 _5413_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4018__B _4283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2680__A2 _2594_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _4954_/A vssd1 vssd1 vccd1 vccd1 _5613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _5564_/Q vssd1 vssd1 vccd1 vccd1 _3905_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2761__B _2761_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5775__D _5775_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _4875_/X _4876_/X _4233_/Y _4877_/X vssd1 vssd1 vccd1 vccd1 _5584_/D sky130_fd_sc_hd__a211o_1
XFILLER_71_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3836_ _4117_/A vssd1 vssd1 vccd1 vccd1 _3836_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4969__A _4990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3767_ _3979_/A vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5506_ _5635_/CLK _5506_/D vssd1 vssd1 vccd1 vccd1 _5506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2718_ _5368_/Q _2613_/X _2717_/Y vssd1 vssd1 vccd1 vccd1 _2787_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__4688__B _4688_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3698_ _3698_/A vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__buf_4
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput330 _3621_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[23] sky130_fd_sc_hd__buf_2
X_5437_ _5446_/CLK _5437_/D vssd1 vssd1 vccd1 vccd1 _5437_/Q sky130_fd_sc_hd__dfxtp_1
X_2649_ _5751_/Q _2577_/X _2648_/Y _2559_/X _2569_/X vssd1 vssd1 vccd1 vccd1 _2650_/B
+ sky130_fd_sc_hd__o2111ai_4
Xoutput341 _3553_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__3145__A0 _5167_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput352 _2942_/X vssd1 vssd1 vccd1 vccd1 ksc_we_o sky130_fd_sc_hd__buf_2
Xoutput363 _3017_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput374 _3039_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[29] sky130_fd_sc_hd__buf_2
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5368_ _5695_/CLK _5368_/D vssd1 vssd1 vccd1 vccd1 _5368_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput385 _5807_/A vssd1 vssd1 vccd1 vccd1 spi_cyc_o sky130_fd_sc_hd__buf_2
XFILLER_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput396 _3172_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[19] sky130_fd_sc_hd__buf_2
XANTENNA__4893__B1 _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4200__C _4252_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_1_0_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _5323_/D sky130_fd_sc_hd__clkbuf_1
X_5299_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5308_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3448__A1 _3267_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5031__C _5039_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2671__B _2695_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5685__D _5685_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3259__S _4803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4581__C1 _4576_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input63_A cpu_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4884__B1 _4872_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output317_A _3578_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3023__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5401__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2662__A2 _2658_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3958__A _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4201__B_N _4076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5595__D _5595_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5551__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3169__S _3192_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4670_ _4778_/C vssd1 vssd1 vccd1 vccd1 _4690_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3621_ _3621_/A vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4167__A2 _4091_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3693__A _5068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3375__A0 _4329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3552_ _3558_/A _3565_/B _4915_/A vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__and3_1
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5116__A1 _5695_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3483_ _3483_/A vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4301__B _4310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5116__B2 _3756_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3127__A0 _5160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5222_/A vssd1 vssd1 vccd1 vccd1 _5740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5153_ _5153_/A vssd1 vssd1 vccd1 vccd1 _5711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4955__C _4955_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _4059_/X _4649_/B _4103_/Y _4007_/X vssd1 vssd1 vccd1 vccd1 _4104_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4627__B1 _3821_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4035_ _5783_/Q _3915_/X _4026_/X _4034_/Y vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__o22ai_4
XFILLER_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2653__A2 _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2772__A _4117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5052__B1 _3540_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4690__C _4690_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4937_ _4937_/A vssd1 vssd1 vccd1 vccd1 _5607_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3079__S _3102_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4868_ _4064_/X _4065_/X _4856_/X _4857_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _5573_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4699__A _4699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3819_ _4253_/D vssd1 vssd1 vccd1 vccd1 _4043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _5540_/Q _4780_/X _4798_/X _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _5540_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5107__A1 _5099_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4211__B _5304_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4866__B1 _4856_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput182 _4010_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_88_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput193 _4168_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[22] sky130_fd_sc_hd__buf_2
XANTENNA__2947__A _3144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5424__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4881__A3 _4847_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2892__A2 _2882_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2644__A2 _5261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3841__A1 _3813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2682__A _5373_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4402__A _4439_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5217__B _5225_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3873__A_N _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output267_A _3443_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3109__A0 _5152_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3018__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2576__B _2616_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2883__A2 _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4085__A1 _3977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3688__A _3742_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2592__A input7/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _5800_/CLK _5771_/D vssd1 vssd1 vccd1 vccd1 _5771_/Q sky130_fd_sc_hd__dfxtp_1
X_2983_ _5741_/Q input30/X _3233_/S vssd1 vssd1 vccd1 vccd1 _5223_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3200__B _3221_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4722_ _4722_/A _4731_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__and3_1
X_4653_ _5474_/Q _4652_/X _4145_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _5474_/D sky130_fd_sc_hd__a211o_1
XFILLER_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput40 cpu_dat_i[14] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
X_3604_ _4289_/D vssd1 vssd1 vccd1 vccd1 _3633_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4312__A _4322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput51 cpu_dat_i[24] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
X_4584_ _4617_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__clkbuf_2
Xinput62 cpu_dat_i[5] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 gpio_ack_i vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__buf_4
XFILLER_50_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3899__B2 _3808_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput84 gpio_dat_i[19] vssd1 vssd1 vccd1 vccd1 _4116_/C sky130_fd_sc_hd__clkbuf_1
Xinput95 gpio_dat_i[29] vssd1 vssd1 vccd1 vccd1 _4257_/C sky130_fd_sc_hd__clkbuf_1
X_3535_ _4304_/B _5595_/Q _3564_/S vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3891__B_N _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2571__A1 _5361_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5447__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3466_ _3654_/S vssd1 vssd1 vccd1 vccd1 _3652_/S sky130_fd_sc_hd__buf_2
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5205_ _5223_/A _5215_/B _5205_/C vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__or3_1
XANTENNA__2767__A _2795_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3397_ _3412_/A _3397_/B _4724_/C vssd1 vssd1 vccd1 vccd1 _3398_/A sky130_fd_sc_hd__and3_1
XFILLER_83_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5143__A _5152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5136_ _5136_/A _5154_/B _5236_/A vssd1 vssd1 vccd1 vccd1 _5137_/A sky130_fd_sc_hd__and3_1
XANTENNA__5597__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4982__A _4982_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5067_ _4889_/X _5060_/X _5066_/X _5061_/X _3792_/B vssd1 vssd1 vccd1 vccd1 _5663_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_61_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4018_ _4283_/A _4283_/B _4283_/C _4018_/D vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__and4_2
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3598__A _3613_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3587__A0 _4335_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4784__C1 _4783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4579__D _4596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2562__A1 _2675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input165_A spi_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2677__A _5367_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5053__A _5056_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A cpu_adr_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4067__A1 _4059_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5016__B1 _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3301__A _3303_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output384_A _2995_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3447__S _3451_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5228__A _5228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3674__C _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2553__A1 _5360_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3971__A _4265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3320_ _3320_/A vssd1 vssd1 vccd1 vccd1 _3320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _5128_/C _5316_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__mux2_8
XANTENNA__5098__A3 _5090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3182__S _3204_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ _4351_/A _5408_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _4514_/C sky130_fd_sc_hd__mux2_1
XFILLER_80_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2856__A2 _2949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2608__A2 _2549_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4307__A _4307_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3211__A _3211_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4026__B _4026_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__A0 _4324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5754_ _5767_/CLK _5754_/D vssd1 vssd1 vccd1 vccd1 _5754_/Q sky130_fd_sc_hd__dfxtp_1
X_2966_ _4386_/A _5422_/Q _3235_/S vssd1 vssd1 vccd1 vccd1 _4550_/C sky130_fd_sc_hd__mux2_1
XFILLER_91_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4705_ _4724_/A _4714_/B _4705_/C vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__or3_1
XANTENNA__5783__D _5783_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5685_ _5692_/CLK _5685_/D vssd1 vssd1 vccd1 vccd1 _5685_/Q sky130_fd_sc_hd__dfxtp_1
X_2897_ _2925_/A _2925_/B _2911_/B vssd1 vssd1 vccd1 vccd1 _4295_/C sky130_fd_sc_hd__and3_2
XFILLER_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2792__A1 _2610_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5138__A _5152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3584__C _4938_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4042__A _4059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4636_ _4638_/A _4636_/B vssd1 vssd1 vccd1 vccd1 _5461_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4977__A _4977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4567_ _4567_/A vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__buf_8
XFILLER_85_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__B1 _3733_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3518_ _3526_/A _5653_/Q vssd1 vssd1 vccd1 vccd1 _3519_/A sky130_fd_sc_hd__and2_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _4514_/A _4498_/B _4498_/C vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__or3_1
XFILLER_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3449_ _4297_/A _5488_/Q _3453_/S vssd1 vssd1 vccd1 vccd1 _4674_/C sky130_fd_sc_hd__mux2_1
XFILLER_98_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__A2 _2750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3105__B _3105_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2701__D1 _2700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5119_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4049__A1 _3977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5246__B1 _2813_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3272__A2 _3268_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2663__C _2663_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4206__D1 _4117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2960__A _3252_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4221__A1 _4059_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5612__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5693__D _5693_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5048__A _5048_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2783__A1 _2813_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5762__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3791__A _4171_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2838__A2 _2837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5237__B1 _2761_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2854__B _3710_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3799__B1 _5559_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__C _4667_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4127__A _4127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3031__A _3031_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3966__A _4036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2820_ _5762_/Q _2577_/X _2819_/Y _2606_/X vssd1 vssd1 vccd1 vccd1 _2820_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3685__B _5270_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2751_ _5360_/Q vssd1 vssd1 vccd1 vccd1 _2751_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2682_ _5373_/Q vssd1 vssd1 vccd1 vccd1 _2682_/Y sky130_fd_sc_hd__inv_2
X_5470_ _5798_/CLK _5470_/D vssd1 vssd1 vccd1 vccd1 _5470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _4421_/A _4439_/C _2932_/D vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__or3b_1
XANTENNA__4797__A _4797_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _5338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3303_ _3303_/A _5543_/Q vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__and2_1
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4283_ _4283_/A _4283_/B _4283_/C _4283_/D vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__and4_2
XANTENNA__3851__D _3851_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4279__A1 _3763_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2748__C _2782_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3206__A _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _5205_/C _5348_/Q _3234_/S vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__mux2_8
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5124__C _5124_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3183_/A _3165_/B _4508_/A vssd1 vssd1 vccd1 vccd1 _3166_/A sky130_fd_sc_hd__and3_1
XFILLER_80_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4963__C _4963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3096_ _5148_/C _5324_/Q _3132_/S vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__mux2_8
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5778__D _5778_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4037__A _4196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5635__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5806_ _5806_/A vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2780__A _2780_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4203__A1 _5478_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3998_ _3998_/A vssd1 vssd1 vccd1 vccd1 _3998_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5737_ _5737_/CLK _5737_/D vssd1 vssd1 vccd1 vccd1 _5737_/Q sky130_fd_sc_hd__dfxtp_1
X_2949_ _2949_/A vssd1 vssd1 vccd1 vccd1 _3157_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5785__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2765__A1 _2585_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3962__B1 _5567_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _5690_/CLK _5668_/D vssd1 vssd1 vccd1 vccd1 _5668_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _3824_/A _3857_/A _4971_/A vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__o21ai_4
X_5599_ _5641_/CLK _5599_/D vssd1 vssd1 vccd1 vccd1 _5599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4500__A _4500_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2658__C _2695_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A ksc_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2674__B _2779_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5688__D _5688_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__B _5655_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4592__D _4596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3245__A2 _2882_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__A3 _3714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2690__A _5379_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input93_A gpio_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3936__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2756__A1 _2752_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4410__A _5228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5225__B _5225_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3181__A1 _5338_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5508__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output347_A _3649_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3026__A _3026_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4130__B1 _4129_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2865__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5658__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5598__D _5598_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4970_ _4970_/A vssd1 vssd1 vccd1 vccd1 _5620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4433__A1 _5261_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3921_ _3921_/A1 _4528_/A _3714_/X _3920_/Y vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__a31oi_4
XFILLER_75_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3696__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3852_ _4265_/B vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2803_ _2632_/Y _2565_/X _2932_/B vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4304__B _4304_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3783_ _5454_/Q _4444_/A _3782_/X vssd1 vssd1 vccd1 vccd1 _3783_/Y sky130_fd_sc_hd__a21oi_4
X_5522_ _5635_/CLK _5522_/D vssd1 vssd1 vccd1 vccd1 _5522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3944__B1 _3943_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2734_ _2761_/C _2761_/D _2734_/C _2761_/B vssd1 vssd1 vccd1 vccd1 _2736_/B sky130_fd_sc_hd__nand4_4
XFILLER_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5453_ _5695_/CLK _5453_/D vssd1 vssd1 vccd1 vccd1 _5453_/Q sky130_fd_sc_hd__dfxtp_1
X_2665_ _2736_/A _2665_/B _2665_/C vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__nand3_4
XFILLER_86_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3862__C _3862_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4404_ _5361_/Q _4400_/X _2570_/Y _4379_/X vssd1 vssd1 vccd1 vccd1 _5361_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4320__A _4320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5384_ _5731_/CLK _5384_/D vssd1 vssd1 vccd1 vccd1 _5384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2596_ _2707_/A _2592_/Y _2549_/X _2595_/Y _2691_/A vssd1 vssd1 vccd1 vccd1 _2596_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__2759__B _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4335_ _4344_/A _4335_/B vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__and2_1
Xclkbuf_opt_1_0_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_1_CLK/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _2728_/A _3716_/X _5483_/Q vssd1 vssd1 vccd1 vccd1 _4266_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__4974__B _4997_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4121__B1 _4120_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3217_ _3217_/A vssd1 vssd1 vccd1 vccd1 _3217_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2775__A _5802_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4197_ _4197_/A vssd1 vssd1 vccd1 vccd1 _4197_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5151__A _5151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3148_ _3148_/A vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4990__A _4990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _5141_/A _5321_/Q _3102_/S vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__mux2_8
XFILLER_58_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2986__A1 _2973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4214__B _4214_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2738__A1 _2672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__B1 _3933_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3772__C _3772_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4230__A _5584_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4587__D _4596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5800__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2685__A _2761_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5061__A _5102_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__A1 _5484_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2977__A1 _5424_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4405__A _4405_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__B1 _4178_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output297_A _3514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3926__B1 _5565_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5330__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4024__A1_N _3989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4778__C _4778_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5236__A _5236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__A _4140_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2579__B _2616_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4039__A1_N _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4120_ _3940_/X _4046_/X _3975_/X _4119_/Y vssd1 vssd1 vccd1 vccd1 _4120_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5480__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4103__B1 _4101_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _3940_/X _4046_/X _3975_/X _4050_/Y vssd1 vssd1 vccd1 vccd1 _4051_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 cpu_adr_i[12] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
X_3002_ _3002_/A vssd1 vssd1 vccd1 vccd1 _3002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4018__C _4283_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ _4953_/A _4965_/B _4965_/C vssd1 vssd1 vccd1 vccd1 _4954_/A sky130_fd_sc_hd__and3_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3090__A0 _5145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3904_ _5460_/Q _3815_/X _3903_/X vssd1 vssd1 vccd1 vccd1 _3904_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__4315__A _4439_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2761__C _2761_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4884_ _4218_/X _4219_/X _4872_/X _4873_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _5583_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _3832_/X _3833_/X _3835_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _3835_/X sky130_fd_sc_hd__and4bb_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3917__B1 _3916_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3766_ _3766_/A vssd1 vssd1 vccd1 vccd1 _3766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4969__B _4990_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5505_ _5555_/CLK _5505_/D vssd1 vssd1 vccd1 vccd1 _5505_/Q sky130_fd_sc_hd__dfxtp_1
X_2717_ _2715_/Y _2640_/X _2716_/Y _2699_/A _2672_/A vssd1 vssd1 vccd1 vccd1 _2717_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__5791__D _5791_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3697_ _3697_/A _3697_/B _3670_/A1 vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__or3b_4
XANTENNA__4688__C _4688_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5146__A _5146_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5436_ _5446_/CLK _5436_/D vssd1 vssd1 vccd1 vccd1 _5436_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput320 _3589_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[14] sky130_fd_sc_hd__buf_2
X_2648_ input9/X _2761_/B _2761_/C _2761_/D vssd1 vssd1 vccd1 vccd1 _2648_/Y sky130_fd_sc_hd__nand4b_4
Xoutput331 _3625_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput342 _3556_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__3145__A1 _5332_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput353 _2952_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput364 _2962_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__4985__A _4985_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5367_ _5695_/CLK _5367_/D vssd1 vssd1 vccd1 vccd1 _5367_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput375 _2967_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[2] sky130_fd_sc_hd__buf_2
X_2579_ _5261_/A _2616_/A vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__nor2_4
Xoutput386 _3055_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__4893__A1 _4832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4200__D _4664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput397 _3063_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4322_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__and2_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5298_ _5789_/Q _5289_/X _4127_/X _4135_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5789_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4249_ _4263_/A _4249_/B vssd1 vssd1 vccd1 vccd1 _4249_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3448__A2 _3268_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5031__D _5043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2671__C _2695_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5353__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4581__B1 _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3275__S _3451_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5056__A _5056_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input56_A cpu_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4895__A _4947_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4884__A1 _4218_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4884__B2 _4873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3304__A _3304_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3023__B _5442_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output212_A _3285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2662__A3 _2613_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A0 _4310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3620_ _3630_/A _3620_/B _4963_/C vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__and3_1
XFILLER_35_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3375__A1 _5502_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3551_ _4312_/B _5599_/Q _3564_/S vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5116__A2 _2882_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3482_ _3482_/A _5637_/Q vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__and2_1
XANTENNA__3127__A1 _5329_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5221_ _5221_/A _5225_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__and3_1
XFILLER_48_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5152_ _5152_/A _5167_/B _5152_/C vssd1 vssd1 vccd1 vccd1 _5153_/A sky130_fd_sc_hd__or3_1
XFILLER_97_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2886__B1 _2885_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4103_ _3997_/X _4062_/X _4101_/X _4102_/X _4005_/X vssd1 vssd1 vccd1 vccd1 _4103_/Y
+ sky130_fd_sc_hd__o221ai_4
X_5083_ _5075_/X _4890_/X _5070_/X _5076_/X _3970_/B vssd1 vssd1 vccd1 vccd1 _5672_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_42_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4627__A1 _5456_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4088__C1 _3946_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4034_ _3887_/X _4644_/B _4033_/Y _4007_/X vssd1 vssd1 vccd1 vccd1 _4034_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__2638__B1 _2932_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5376__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5786__D _5786_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5052__A1 _5656_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5052__B2 _5034_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4936_ _4936_/A _4940_/B _4940_/C vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__and3_1
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4260__C1 _4259_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2810__B1 _2682_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4867_ _4859_/X _4860_/X _4050_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5572_/D sky130_fd_sc_hd__a211o_1
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3818_ _4076_/A vssd1 vssd1 vccd1 vccd1 _3818_/X sky130_fd_sc_hd__clkbuf_1
X_4798_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4699__B _4714_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3749_ _2859_/Y _3455_/A _5058_/B _3697_/X vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__a211oi_4
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3095__S _3108_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5107__A2 _5094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5419_ _5695_/CLK _5419_/D vssd1 vssd1 vccd1 vccd1 _5419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4866__A1 _4031_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput183 _4022_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__4866__B2 _4857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput194 _4183_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3124__A _3124_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2629__B1 _2628_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5719__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3841__A2 _3822_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input110_A ksc_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5696__D _5696_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2801__B1 _3979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3794__A _4265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5217__C _5231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3109__A1 _5326_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3034__A _3038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2576__C _5261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5399__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3969__A _4171_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4085__A2 _3978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5800_/CLK _5770_/D vssd1 vssd1 vccd1 vccd1 _5770_/Q sky130_fd_sc_hd__dfxtp_1
X_2982_ _2973_/X _2974_/X _4556_/A vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3200__C _4522_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4721_ _4746_/A vssd1 vssd1 vccd1 vccd1 _4741_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4652_ _4652_/A vssd1 vssd1 vccd1 vccd1 _4652_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3603_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3620_/B sky130_fd_sc_hd__clkbuf_1
Xinput30 cpu_adr_i[6] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput41 cpu_dat_i[15] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _5435_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4312__B _4312_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput52 cpu_dat_i[25] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 cpu_dat_i[6] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput74 gpio_dat_i[0] vssd1 vssd1 vccd1 vccd1 _3732_/C sky130_fd_sc_hd__clkbuf_4
Xinput85 gpio_dat_i[1] vssd1 vssd1 vccd1 vccd1 _3772_/C sky130_fd_sc_hd__buf_2
X_3534_ _3654_/S vssd1 vssd1 vccd1 vccd1 _3564_/S sky130_fd_sc_hd__buf_2
Xinput96 gpio_dat_i[2] vssd1 vssd1 vccd1 vccd1 _3797_/C sky130_fd_sc_hd__buf_2
XANTENNA__2571__A2 _2565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3465_ _4289_/D vssd1 vssd1 vccd1 vccd1 _3654_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5204_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5223_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3396_ _4342_/A _5508_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _4724_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2767__B _2795_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5143__B _5143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5135_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5258__D1 _4377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5066_ _5066_/A vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4982__B _4997_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4017_ _4011_/Y _3848_/X _4016_/Y vssd1 vssd1 vccd1 vccd1 _4017_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3598__B _3601_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3587__A1 _5609_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4784__B1 _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4919_ _5005_/B vssd1 vssd1 vccd1 vccd1 _4938_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4503__A _4514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3119__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2562__A2 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input158_A spi_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5053__B _5657_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5541__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4067__A2 _4647_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3275__A0 _4396_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A cpu_adr_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5691__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5016__A1 _5638_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5016__B2 _5011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3301__B _5542_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4116__C _4116_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__C1 _2540_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output377_A _3043_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3029__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2553__A2 _2540_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3463__S _3645_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3250_ _5701_/Q input70/X _3250_/S vssd1 vssd1 vccd1 vccd1 _5128_/C sky130_fd_sc_hd__mux2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3181_ _5181_/C _5338_/Q _3192_/S vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__mux2_8
XFILLER_67_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2710__C1 _2606_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3266__B1 _4769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4026__C _4159_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__A1 _5604_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5753_ _5767_/CLK _5753_/D vssd1 vssd1 vccd1 vccd1 _5753_/Q sky130_fd_sc_hd__dfxtp_1
X_2965_ _5215_/C _5352_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__mux2_8
XFILLER_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4704_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4323__A _4323_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5684_ _5690_/CLK _5684_/D vssd1 vssd1 vccd1 vccd1 _5684_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5414__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2896_ _2909_/A _2909_/B _2909_/C _2929_/B vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__and4_1
XANTENNA__5138__B _5143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2792__A2 _5227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4635_ _5460_/Q _4623_/X _3903_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _5460_/D sky130_fd_sc_hd__a211o_1
XFILLER_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4566_ _5428_/Q _4563_/X _5807_/A _4564_/X _4565_/X vssd1 vssd1 vccd1 vccd1 _5428_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3741__A1 _3720_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3517_ _3517_/A vssd1 vssd1 vccd1 vccd1 _3526_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3741__B2 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2778__A _4098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4497_ _4497_/A vssd1 vssd1 vccd1 vccd1 _5401_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5154__A _5154_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3448_ _3267_/X _3268_/X _4671_/A vssd1 vssd1 vccd1 vccd1 _3448_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4993__A _4993_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _4331_/B _5503_/Q _3400_/S vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__mux2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2701__C1 _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3105__C _4481_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5697_/Q _2927_/A _5060_/X _5114_/X _4848_/X vssd1 vssd1 vccd1 vccd1 _5697_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4049__A2 _3978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5246__A1 _5752_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5654_/Q _5033_/X _3540_/A _5034_/X _5045_/X vssd1 vssd1 vccd1 vccd1 _5654_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3402__A _3402_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__D _2761_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4206__C1 _4205_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4221__A2 _4658_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2783__A2 _2848_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5064__A _5064_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5237__A1 _5746_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3248__A0 _4299_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4408__A _4600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__A1 _4830_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4127__B _4127_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__D _4665_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5437__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3966__B _3966_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3685__C _3685_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2750_ _2750_/A vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4143__A _4252_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2681_ _2813_/A _2615_/X _2680_/Y _2574_/A vssd1 vssd1 vccd1 vccd1 _4417_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__5587__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4420_ _5369_/Q _5238_/A _2721_/Y _4299_/A vssd1 vssd1 vccd1 vccd1 _5369_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2598__A _2647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4351_ _4351_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__or2_1
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3193__S _3204_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3302_ _3302_/A vssd1 vssd1 vccd1 vccd1 _3302_/X sky130_fd_sc_hd__clkbuf_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _4276_/Y _3848_/X _4281_/Y vssd1 vssd1 vccd1 vccd1 _4282_/Y sky130_fd_sc_hd__o21ai_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4279__A2 _3766_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2748__D _2935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _5733_/Q input59/X _3233_/S vssd1 vssd1 vccd1 vccd1 _5205_/C sky130_fd_sc_hd__mux2_2
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _4344_/B _5405_/Q _3209_/S vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3239__A0 _5120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4318__A _4322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3095_ _5709_/Q input64/X _3108_/S vssd1 vssd1 vccd1 vccd1 _5148_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3222__A _3222_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5805_ _5805_/A vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2780__B _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5794__D _5794_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3368__S _3396_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3997_ _4147_/A vssd1 vssd1 vccd1 vccd1 _3997_/X sky130_fd_sc_hd__buf_4
XANTENNA__4203__A2 _4074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5149__A _5149_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3411__A0 _4351_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5736_ _5765_/CLK _5736_/D vssd1 vssd1 vccd1 vccd1 _5736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2948_ _5210_/C _5350_/Q _3234_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__mux2_8
XANTENNA__2765__A2 _2790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3962__A1 _3961_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5667_ _5802_/CLK _5667_/D vssd1 vssd1 vccd1 vccd1 _5667_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4988__A _4988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2879_ _2879_/A vssd1 vssd1 vccd1 vccd1 _2925_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4618_ _4618_/A vssd1 vssd1 vccd1 vccd1 _5452_/D sky130_fd_sc_hd__clkbuf_1
X_5598_ _5641_/CLK _5598_/D vssd1 vssd1 vccd1 vccd1 _5598_/Q sky130_fd_sc_hd__dfxtp_1
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _5421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4500__B _4500_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__D _2695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3478__B1 _5007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4228__A _4254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2674__C _2779_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__C _5056_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3650__A0 _4297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5059__A _5059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input86_A gpio_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2756__A2 _2552_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4898__A _4898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3307__A _3307_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5225__C _5231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output242_A _3282_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4130__A1 _4130_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2865__B _2917_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4138__A _4138_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3042__A _3042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4433__A2 input20/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5091__C1 _4041_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3977__A _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3920_ _3794_/X _3919_/X _5461_/Q vssd1 vssd1 vccd1 vccd1 _3920_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__2881__A _4295_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3968__A2_N _5672_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3851_ _4254_/A _4265_/B _4283_/C _3851_/D vssd1 vssd1 vccd1 vccd1 _3851_/X sky130_fd_sc_hd__and4_2
XANTENNA__3188__S _3209_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2802_ _2778_/Y _3403_/A _3961_/A vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__a21oi_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _3878_/A _4283_/B _4283_/C _3782_/D vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__and4_2
X_5521_ _5555_/CLK _5521_/D vssd1 vssd1 vccd1 vccd1 _5521_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3944__A1 _3941_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2733_ _4415_/A _4415_/B _2780_/B _2787_/A _2787_/B vssd1 vssd1 vccd1 vccd1 _2741_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4601__A _4611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5452_ _5586_/CLK _5452_/D vssd1 vssd1 vccd1 vccd1 _5452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2664_ _2593_/X _2594_/X _5756_/Q vssd1 vssd1 vccd1 vccd1 _2665_/C sky130_fd_sc_hd__o21ai_2
XFILLER_86_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4403_ _2752_/Y _2552_/Y _4402_/X vssd1 vssd1 vccd1 vccd1 _5360_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5383_ _5435_/CLK _5383_/D vssd1 vssd1 vccd1 vccd1 _5383_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3862__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4320__B _4333_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2595_ _2593_/X _2594_/X _5749_/Q vssd1 vssd1 vccd1 vccd1 _2595_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3217__A _3217_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2759__C _2759_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2904__C1 _2779_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4334_ _4334_/A vssd1 vssd1 vccd1 vccd1 _5330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4265_ _4265_/A _4265_/B _4265_/C _4265_/D vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__and4_2
XANTENNA__4974__C _4997_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4657__C1 _4621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__A1 _4042_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ _3236_/A _3221_/B _4529_/C vssd1 vssd1 vccd1 vccd1 _3217_/A sky130_fd_sc_hd__and3_1
XANTENNA__5602__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5789__D _5789_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4196_ _4196_/A vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__buf_8
XFILLER_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3147_ _3152_/A _3165_/B _4498_/C vssd1 vssd1 vccd1 vccd1 _3148_/A sky130_fd_sc_hd__and3_1
XFILLER_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3880__B1 _5289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3078_ _5706_/Q input61/X _3126_/S vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4990__B _4990_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5082__C1 _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3887__A _4059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5752__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2986__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3098__S _3146_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4214__C _4240_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2738__A2 _2699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5741_/CLK _5719_/D vssd1 vssd1 vccd1 vccd1 _5719_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3935__B2 _3934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4511__A _4511_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3772__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3561__S _3642_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4648__C1 _4645_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input140_A ksc_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5699__D _5699_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4663__A2 _4542_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3871__B1 _3846_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__C1 _5111_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3623__A0 _4357_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4405__B _4425_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__A1 _4176_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3926__A1 _4830_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output192_A _4156_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4421__A _4421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3037__A _3037_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4887__C1 _4877_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5625__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2876__A _3042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3471__S _3645_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4103__A1 _3997_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4103__B2 _4102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4050_ _4047_/Y _3906_/X _4049_/Y vssd1 vssd1 vccd1 vccd1 _4050_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3001_ _3005_/A _5432_/Q vssd1 vssd1 vccd1 vccd1 _3002_/A sky130_fd_sc_hd__and2_1
Xinput6 cpu_adr_i[13] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5775__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5402__D _5402_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4018__D _4018_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4952_ _4952_/A vssd1 vssd1 vccd1 vccd1 _5612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3500__A _3504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3924__A_N _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3903_ _4283_/A _4079_/B _3903_/C vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__and3_1
XANTENNA__3090__A1 _5323_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4883_ _5235_/A vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__buf_4
XANTENNA__2761__D _2761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3834_ _4099_/A vssd1 vssd1 vccd1 vccd1 _4269_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3917__B2 _3700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3765_ _4257_/D vssd1 vssd1 vccd1 vccd1 _3766_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4969__C _4969_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5504_ _5538_/CLK _5504_/D vssd1 vssd1 vccd1 vccd1 _5504_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3873__C _3873_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2716_ _2607_/A _2549_/A _5753_/Q vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__4331__A _4344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__inv_2
X_5435_ _5435_/CLK _5435_/D vssd1 vssd1 vccd1 vccd1 _5435_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput310 _3476_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[6] sky130_fd_sc_hd__buf_2
X_2647_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2761_/C sky130_fd_sc_hd__clkbuf_4
Xoutput321 _3592_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput332 _3628_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4878__C1 _4877_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput343 _3559_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput354 _2998_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[10] sky130_fd_sc_hd__buf_2
X_5366_ _5695_/CLK _5366_/D vssd1 vssd1 vccd1 vccd1 _5366_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput365 _3020_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[20] sky130_fd_sc_hd__buf_2
XFILLER_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2578_ input6/X vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__inv_2
Xoutput376 _3041_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[30] sky130_fd_sc_hd__buf_2
Xoutput387 _3118_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[10] sky130_fd_sc_hd__buf_2
XANTENNA__4893__A2 _4833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _5322_/D sky130_fd_sc_hd__clkbuf_1
Xoutput398 _3178_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_87_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5297_ _5297_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5788_/D sky130_fd_sc_hd__nand2_1
XFILLER_82_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5162__A _5176_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4248_ _5797_/Q _4091_/X _4240_/X _4247_/Y vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__o22ai_4
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _4176_/Y _4115_/X _4178_/Y vssd1 vssd1 vccd1 vccd1 _4179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5055__C1 _5045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3605__A0 _4346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4506__A _4971_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__A _3410_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3942__B_N _3833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2671__D _2695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4581__A1 _5434_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4581__B2 _4564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5648__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5056__B _5659_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4869__C1 _4861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4884__A2 _4219_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2696__A _2696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5798__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input49_A cpu_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5072__A _5072_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4097__B1 _4096_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5294__C1 _5285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5046__C1 _5045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output205_A _3869_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4416__A _4416_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A1 _5390_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4021__B1 _4017_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3550_ _4988_/B vssd1 vssd1 vccd1 vccd1 _3565_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _3481_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3990__A _3990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5220_ _5220_/A vssd1 vssd1 vccd1 vccd1 _5739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5151_ _5151_/A vssd1 vssd1 vccd1 vccd1 _5710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2886__A1 _2946_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _3961_/X _4003_/X _5575_/Q vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5082_ _5081_/X _5078_/X _5066_/X _5061_/X _3953_/B vssd1 vssd1 vccd1 vccd1 _5671_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4088__B1 _4087_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__A2 _4623_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4033_ _3997_/X _3890_/X _4031_/X _4032_/X _4005_/X vssd1 vssd1 vccd1 vccd1 _4033_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2638__A1 _2632_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4326__A _4441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5052__A2 _5021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _4935_/A vssd1 vssd1 vccd1 vccd1 _5606_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4260__B1 _3758_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2810__A1 _2809_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4866_ _4031_/X _4032_/X _4856_/X _4857_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _5571_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3817_ _4075_/A vssd1 vssd1 vccd1 vccd1 _3817_/X sky130_fd_sc_hd__clkbuf_1
X_4797_ _4797_/A vssd1 vssd1 vccd1 vccd1 _5539_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4699__C _4699_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5157__A _5176_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3748_ _3989_/A vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__buf_4
XANTENNA__4996__A _4996_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_1_0_1_CLK_A clkbuf_1_0_1_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5107__A3 _5066_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3679_ _3979_/A _4746_/A _3678_/X vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__a21oi_1
XFILLER_97_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5418_ _5586_/CLK _5418_/D vssd1 vssd1 vccd1 vccd1 _5418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4866__A2 _4032_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput184 _4036_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[14] sky130_fd_sc_hd__buf_2
X_5349_ _5767_/CLK _5349_/D vssd1 vssd1 vccd1 vccd1 _5349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput195 _4195_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3405__A _3412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5276__C1 _5310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2629__A1 _5358_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5320__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input103_A gpio_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4251__B1 _4250_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2801__A1 _3980_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5470__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2868__A1 _3670_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3315__A _3315_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3034__B _5447_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output322_A _3595_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5019__C1 _4823_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _4392_/B _5425_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__mux2_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4242__B1 _4241_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4720_ _4720_/A vssd1 vssd1 vccd1 vccd1 _5506_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4651_ _4651_/A _4651_/B vssd1 vssd1 vccd1 vccd1 _5473_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3602_ _3602_/A vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__clkbuf_1
Xinput20 cpu_adr_i[26] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_4
Xinput31 cpu_adr_i[7] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _4592_/A _5435_/Q _4665_/D _4596_/D vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__and4_1
XFILLER_50_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 cpu_dat_i[16] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_0_CLK_A CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput53 cpu_dat_i[26] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 cpu_dat_i[7] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
Xinput75 gpio_dat_i[10] vssd1 vssd1 vccd1 vccd1 _3959_/C sky130_fd_sc_hd__buf_2
X_3533_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__clkbuf_4
Xinput86 gpio_dat_i[20] vssd1 vssd1 vccd1 vccd1 _4131_/C sky130_fd_sc_hd__clkbuf_2
Xinput97 gpio_dat_i[30] vssd1 vssd1 vccd1 vccd1 _4269_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3464_ _2924_/X _2927_/X _4995_/C vssd1 vssd1 vccd1 vccd1 _3464_/X sky130_fd_sc_hd__o21a_1
X_5203_ _5203_/A vssd1 vssd1 vccd1 vccd1 _5732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3395_ _3431_/A vssd1 vssd1 vccd1 vccd1 _3412_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5134_/A vssd1 vssd1 vccd1 vccd1 _5703_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5143__C _5143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5258__C1 _5228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5343__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5065_ _5662_/Q _4988_/A _3750_/X _5065_/B2 _5111_/B vssd1 vssd1 vccd1 vccd1 _5662_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4982__C _4997_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4016_ _4628_/A _3857_/X _5099_/A _4015_/Y vssd1 vssd1 vccd1 vccd1 _4016_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5797__D _5797_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3598__C _4951_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5493__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4233__B1 _4232_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4784__A1 _5532_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _4968_/A vssd1 vssd1 vccd1 vccd1 _5005_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4784__B2 _4782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4503__B _4524_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4849_ _3662_/Y _3678_/X _4847_/X _3864_/Y _4848_/X vssd1 vssd1 vccd1 vccd1 _5561_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3744__C1 _3743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3135__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5053__C _5056_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5249__C1 _5238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2974__A _4295_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3275__A1 _5531_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5500__D _5500_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5016__A2 _5010_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4116__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2786__B1 _2658_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output272_A _3358_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5366__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3045__A _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3180_ _5723_/Q input48/X _3223_/S vssd1 vssd1 vccd1 vccd1 _5181_/C sky130_fd_sc_hd__mux2_2
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2710__B1 _2709_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3699__B _3699_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3266__A1 _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5410__D _5410_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4026__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4604__A _4611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5752_ _5767_/CLK _5752_/D vssd1 vssd1 vccd1 vccd1 _5752_/Q sky130_fd_sc_hd__dfxtp_1
X_2964_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3251_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4703_ _5270_/A vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__buf_2
X_2895_ _3329_/A vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5683_ _5690_/CLK _5683_/D vssd1 vssd1 vccd1 vccd1 _5683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5138__C _5138_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4634_ _4638_/A _4634_/B vssd1 vssd1 vccd1 vccd1 _5459_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4565_ _4891_/A vssd1 vssd1 vccd1 vccd1 _4565_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5709__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3654__S _3654_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3516_ _3516_/A vssd1 vssd1 vccd1 vccd1 _3516_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3741__A2 _3722_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4496_ _4496_/A _4500_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__and3_1
XFILLER_85_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5154__B _5154_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3447_ _4292_/B _5487_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3431_/A vssd1 vssd1 vccd1 vccd1 _3393_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2701__B1 _2698_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__A _2794_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5117_ _5696_/Q _2899_/A _5070_/X _4847_/X _4848_/X vssd1 vssd1 vccd1 vccd1 _5696_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5170__A _5170_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5246__A2 _5234_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5320__D _5320_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4217__C _4217_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4206__B1 _3768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4514__A _4514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2783__A3 _2848_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5389__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3564__S _3564_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3193__A0 _4355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input170_A spi_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4189__B_N _3861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input31_A cpu_adr_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5237__A2 _5234_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3248__A1 _5385_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3312__B _5547_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__A2 _3737_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4127__C _4159_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4424__A _4424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4143__B _4143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2680_ _2593_/X _2594_/X _5752_/Q vssd1 vssd1 vccd1 vccd1 _2680_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2879__A _2879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5255__A _5255_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4350_ _4350_/A vssd1 vssd1 vccd1 vccd1 _5337_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2598__B _2686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3301_ _3303_/A _5542_/Q vssd1 vssd1 vccd1 vccd1 _3302_/A sky130_fd_sc_hd__and2_1
XANTENNA__2931__B1 _5372_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4281_ _4628_/A _3857_/X _5099_/A _4280_/Y vssd1 vssd1 vccd1 vccd1 _4281_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5405__D _5405_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3232_/X sky130_fd_sc_hd__clkbuf_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3163_ _3163_/A vssd1 vssd1 vccd1 vccd1 _3209_/S sky130_fd_sc_hd__buf_2
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3503__A _3503_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _4617_/A vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3239__A1 _5313_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4318__B _4318_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4436__B1 _4402_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4334__A _4334_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2780__C _2780_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3996_ _3996_/A1 _3954_/X _3994_/X _3995_/Y vssd1 vssd1 vccd1 vccd1 _4642_/B sky130_fd_sc_hd__a31oi_4
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3947__C1 _3946_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5735_ _5737_/CLK _5735_/D vssd1 vssd1 vccd1 vccd1 _5735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3234_/S sky130_fd_sc_hd__buf_4
XANTENNA__3411__A1 _5512_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5531__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3962__A2 _3737_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5666_ _5694_/CLK _5666_/D vssd1 vssd1 vccd1 vccd1 _5666_/Q sky130_fd_sc_hd__dfxtp_1
X_2878_ _2878_/A _2917_/A vssd1 vssd1 vccd1 vccd1 _2887_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4988__B _4988_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4617_ _4617_/A _4617_/B _4796_/C vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__and3_1
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5597_ _5641_/CLK _5597_/D vssd1 vssd1 vccd1 vccd1 _5597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3175__A0 _5178_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5165__A _5165_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4548_ _4548_/A _4556_/B _4569_/A vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__and3_1
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5681__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4500__C _4512_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5315__D _5315_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4479_ _4479_/A vssd1 vssd1 vccd1 vccd1 _5394_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3478__A1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4509__A _4509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__A _3413_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4228__B _4228_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2674__D _2935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__D _5056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__A0 _4396_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3650__A1 _5592_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4898__B _4915_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input79_A gpio_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2699__A _2699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5075__A _5096_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4130__A2 _4449_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output235_A _3330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3323__A _3325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3874__D1 _3331_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5404__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3042__B _5451_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output402_A _3201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5091__B1 _5076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4433__A3 _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5554__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _3850_/A vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2801_ _3980_/A _3977_/A _3979_/A vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__o21ai_4
X_3781_ _4265_/C vssd1 vssd1 vccd1 vccd1 _4283_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3993__A _4127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5635_/CLK _5520_/D vssd1 vssd1 vccd1 vccd1 _5520_/Q sky130_fd_sc_hd__dfxtp_1
X_2732_ _5367_/Q _2621_/X _4417_/B vssd1 vssd1 vccd1 vccd1 _2780_/B sky130_fd_sc_hd__o21ai_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3944__A2 _3906_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5451_ _5531_/CLK _5451_/D vssd1 vssd1 vccd1 vccd1 _5451_/Q sky130_fd_sc_hd__dfxtp_1
X_2663_ _2761_/C _2761_/D _2663_/C _2761_/B vssd1 vssd1 vccd1 vccd1 _2665_/B sky130_fd_sc_hd__nand4_4
XANTENNA__4601__B _5443_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4402_ _4439_/C vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2594_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__clkbuf_4
X_5382_ _5800_/CLK _5382_/D vssd1 vssd1 vccd1 vccd1 _5382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2904__B1 _2814_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2759__D _2864_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4333_ _4333_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__or2_1
XFILLER_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4264_ _5691_/Q _4986_/A _3846_/A _4264_/B2 vssd1 vssd1 vccd1 vccd1 _5111_/A sky130_fd_sc_hd__a22oi_4
XANTENNA__4657__B1 _4202_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3215_ _4364_/A _5414_/Q _3235_/S vssd1 vssd1 vccd1 vccd1 _4529_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4121__A2 _4113_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4329__A _4329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4195_ _4195_/A _4195_/B vssd1 vssd1 vccd1 vccd1 _4195_/Y sky130_fd_sc_hd__nor2_8
XFILLER_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3146_ _4338_/A _5402_/Q _3146_/S vssd1 vssd1 vccd1 vccd1 _4498_/C sky130_fd_sc_hd__mux2_1
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3880__A1 _3707_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3077_ _3250_/S vssd1 vssd1 vccd1 vccd1 _3126_/S sky130_fd_sc_hd__buf_2
XANTENNA__4990__C _4990_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5082__B1 _5061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3379__S _3400_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4999__A _5128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3396__A0 _4342_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3979_ _3979_/A vssd1 vssd1 vccd1 vccd1 _3979_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4214__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5718_ _5765_/CLK _5718_/D vssd1 vssd1 vccd1 vccd1 _5718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5649_ _5659_/CLK _5649_/D vssd1 vssd1 vccd1 vccd1 _5649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5427__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4648__B1 _4079_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4227__B_N _4076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input133_A ksc_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3871__A1 _5666_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5577__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3871__B2 _5073_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__B1 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A1 _5619_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__A2 _4115_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4702__A _4702_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3926__A2 _3737_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output185_A _4054_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4421__B _4439_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3139__A0 _5165_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3318__A _3318_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4887__B1 _4259_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output352_A _2942_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4103__A2 _4062_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3000_ _3000_/A vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 cpu_adr_i[14] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3988__A _5068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4951_ _4963_/A _4963_/B _4951_/C vssd1 vssd1 vccd1 vccd1 _4952_/A sky130_fd_sc_hd__or3_1
XANTENNA__3199__S _3209_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3500__B _5645_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3902_ _3817_/X _3818_/X _3902_/C _4043_/D vssd1 vssd1 vccd1 vccd1 _3903_/C sky130_fd_sc_hd__and4bb_1
XFILLER_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _4875_/X _4876_/X _4207_/Y _4877_/X vssd1 vssd1 vccd1 vccd1 _5582_/D sky130_fd_sc_hd__a211o_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3833_ _4083_/A vssd1 vssd1 vccd1 vccd1 _3833_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4612__A _4612_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3764_ _3980_/A vssd1 vssd1 vccd1 vccd1 _4257_/D sky130_fd_sc_hd__clkbuf_2
X_5503_ _5538_/CLK _5503_/D vssd1 vssd1 vccd1 vccd1 _5503_/Q sky130_fd_sc_hd__dfxtp_1
X_2715_ _2715_/A vssd1 vssd1 vccd1 vccd1 _2715_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3873__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4331__B _4331_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3695_ _3989_/A vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput300 _3521_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[26] sky130_fd_sc_hd__buf_2
X_5434_ _5435_/CLK _5434_/D vssd1 vssd1 vccd1 vccd1 _5434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2646_ _2809_/A _2750_/A _5366_/Q vssd1 vssd1 vccd1 vccd1 _2650_/A sky130_fd_sc_hd__o21ai_1
Xoutput311 _3478_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[7] sky130_fd_sc_hd__buf_2
Xoutput322 _3595_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__4878__B1 _4151_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput333 _3631_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_47_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput344 _3563_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput355 _3000_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[11] sky130_fd_sc_hd__buf_2
X_2577_ _2785_/A vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__clkbuf_4
X_5365_ _5765_/CLK _5365_/D vssd1 vssd1 vccd1 vccd1 _5365_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput366 _3022_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput377 _3043_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[31] sky130_fd_sc_hd__buf_2
XFILLER_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput388 _3124_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4316_ _4316_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__or2_1
XFILLER_82_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput399 _3184_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[21] sky130_fd_sc_hd__buf_2
X_5296_ _5787_/Q _5289_/X _4094_/X _4104_/Y _5285_/X vssd1 vssd1 vccd1 vccd1 _5787_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5162__B _5167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4247_ _3813_/X _4660_/B _4246_/Y _3840_/X vssd1 vssd1 vccd1 vccd1 _4247_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4059__A _4059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4178_ _3763_/A _3766_/A _3768_/A _4177_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4178_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3853__A1 _2728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3898__A _3898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3129_ _3152_/A _3134_/B _4491_/A vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__and3_1
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5055__B1 _3540_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3605__A1 _5614_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4566__C1 _4565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4522__A _4522_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3952__A2_N _5671_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4581__A2 _4563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5056__C _5056_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4869__B1 _4086_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2696__B _2696_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5072__B _5111_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5503__D _5503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__A1 _4097_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5294__B1 _4058_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5046__B1 _5029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3601__A _3613_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4432__A _4432_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__A1 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__B2 _4020_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3480_ _3482_/A _5636_/Q vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__and2_1
XFILLER_13_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2887__A _2909_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5742__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5150_ _5150_/A _5154_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__and3_1
XANTENNA__3795__B1_N _5455_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2886__A2 _5208_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4101_ _4098_/X _3958_/X _3998_/X _4100_/X vssd1 vssd1 vccd1 vccd1 _4101_/X sky130_fd_sc_hd__o211a_1
X_5081_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5413__D _5413_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4088__A1 _4042_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4032_ _3961_/X _4003_/X _5571_/Q vssd1 vssd1 vccd1 vccd1 _4032_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__A2 _2613_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4607__A _5042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3511__A _3515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4934_ _4938_/A _4938_/B _4934_/C vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__or3_1
XANTENNA__4260__A1 _4147_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _5235_/A vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2810__A2 _2750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4342__A _4342_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3816_ _3849_/A vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__clkbuf_1
X_4796_ _4801_/A _5539_/Q _4796_/C vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__and3_1
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5157__B _5167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3747_ _4091_/A vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__buf_6
XFILLER_88_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3678_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5417_ _5531_/CLK _5417_/D vssd1 vssd1 vccd1 vccd1 _5417_/Q sky130_fd_sc_hd__dfxtp_1
X_2629_ _5358_/Q _2621_/X _2628_/Y vssd1 vssd1 vccd1 vccd1 _2864_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__2797__A _2853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__S _3400_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5173__A _5173_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5348_ _5482_/CLK _5348_/D vssd1 vssd1 vccd1 vccd1 _5348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput185 _4054_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput196 _4211_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[25] sky130_fd_sc_hd__buf_2
XANTENNA__3405__B _3416_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5323__D _5323_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5279_ _5773_/Q _5114_/X _5069_/X _3867_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5773_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5276__B1 _3792_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2629__A2 _2621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4517__A _4517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3421__A _3421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5615__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4251__B2 _4141_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2801__A2 _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4252__A _4252_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5765__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input61_A cpu_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2868__A2 _2867_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output315_A _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4427__A _4431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5019__B1 _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3331__A _3331_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _5221_/A _5355_/Q _3229_/S vssd1 vssd1 vccd1 vccd1 _4392_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4242__A1 _4242_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3477__S _3652_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _5472_/Q _4639_/X _4112_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _5472_/D sky130_fd_sc_hd__a211o_1
X_3601_ _3613_/A _3601_/B _4953_/A vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__and3_1
Xinput10 cpu_adr_i[17] vssd1 vssd1 vccd1 vccd1 _2679_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 cpu_adr_i[27] vssd1 vssd1 vccd1 vccd1 _2651_/A sky130_fd_sc_hd__clkbuf_2
X_4581_ _5434_/Q _4563_/X _5807_/A _4564_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _5434_/D
+ sky130_fd_sc_hd__a221o_1
Xinput32 cpu_adr_i[8] vssd1 vssd1 vccd1 vccd1 _2836_/A sky130_fd_sc_hd__buf_6
XANTENNA__5408__D _5408_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput43 cpu_dat_i[17] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 cpu_dat_i[27] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3532_ _3699_/B vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__clkbuf_2
Xinput65 cpu_dat_i[8] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 gpio_dat_i[11] vssd1 vssd1 vccd1 vccd1 _3981_/C sky130_fd_sc_hd__clkbuf_1
Xinput87 gpio_dat_i[21] vssd1 vssd1 vccd1 vccd1 _4149_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput98 gpio_dat_i[31] vssd1 vssd1 vccd1 vccd1 _4278_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3463_ _4386_/A _5630_/Q _3645_/S vssd1 vssd1 vccd1 vccd1 _4995_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3506__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5202_ _5202_/A _5202_/B _5208_/C vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__and3_1
X_3394_ _3394_/A vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5133_ _5152_/A _5143_/B _5133_/C vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__or3_1
XANTENNA__5258__B1 _2819_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4015_ _4012_/Y _4743_/A _4014_/Y vssd1 vssd1 vccd1 vccd1 _4015_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__4337__A _4385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5638__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4233__A1 _4230_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4784__A2 _4780_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5788__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5168__A _5168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3992__B1 _3990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4848_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__buf_4
XANTENNA__4503__C _4503_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4779_ _4779_/A vssd1 vssd1 vccd1 vccd1 _5531_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5318__D _5318_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3744__B1 _3741_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4800__A _5207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3937__A_N _3817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3416__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5053__D _5056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5249__B1 _4891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5078__A _5094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2786__A1 _5759_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3983__B1 _3982_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5806__A _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4710__A _4710_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output265_A _3440_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3326__A _3326_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5589_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2710__A1 _5261_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4157__A _4157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3699__C _5034_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__A2 _2899_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4215__A1 _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5751_ _5767_/CLK _5751_/D vssd1 vssd1 vccd1 vccd1 _5751_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4604__B _5445_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2963_ _5737_/Q input24/X _3233_/S vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__mux2_1
XFILLER_91_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4702_ _4702_/A vssd1 vssd1 vccd1 vccd1 _5499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3974__B1 _3973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5682_ _5692_/CLK _5682_/D vssd1 vssd1 vccd1 vccd1 _5682_/Q sky130_fd_sc_hd__dfxtp_1
X_2894_ _3277_/A vssd1 vssd1 vccd1 vccd1 _3329_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _5458_/Q _4623_/X _3878_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _5458_/D sky130_fd_sc_hd__a211o_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4620__A _4645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4564_ _4590_/A vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__buf_2
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2934__D1 _2779_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3515_ _3515_/A _5652_/Q vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__and2_1
XFILLER_89_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ _4495_/A vssd1 vssd1 vccd1 vccd1 _5400_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3236__A _3236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5154__C _5160_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3446_ _3446_/A vssd1 vssd1 vccd1 vccd1 _3446_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4151__B1 _4150_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3377_ _3377_/A vssd1 vssd1 vccd1 vccd1 _3377_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2701__A1 _5764_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5116_ _5695_/Q _2882_/A _4667_/C _3756_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _5695_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5460__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__B _2852_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5100__C1 _4127_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5047_ _5056_/A _5653_/Q _5056_/C _5056_/D vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__and4_1
XFILLER_61_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5601__D _5601_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__A1 _3763_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4514__B _4524_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3965__B1 _3953_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4530__A _4530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3193__A1 _5410_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input163_A spi_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4142__B1 _4140_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3580__S _3600_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A cpu_adr_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5511__D _5511_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4127__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4705__A _4724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5741_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3956__B1 _3955_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4143__C _4143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output382_A _2990_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5333__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4440__A _4440_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5255__B _5266_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2598__C input8/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3056__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3300_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2931__A1 _5266_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5483__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4280_ _4277_/Y _3828_/X _4279_/Y vssd1 vssd1 vccd1 vccd1 _4280_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4133__B1 _5577_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2895__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3231_ _3236_/A _4542_/B _4536_/A vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__and3_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5271__A _5299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3162_ _5174_/A _5335_/Q _3162_/S vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__mux2_8
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3892__C1 _3891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3093_ _3093_/A vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5421__D _5421_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4436__A1 _2817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4615__A _4615_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3995_ _3794_/X _3919_/X _5465_/Q vssd1 vssd1 vccd1 vccd1 _3995_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__2780__D _2780_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3947__B1 _3945_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5734_ _5765_/CLK _5734_/D vssd1 vssd1 vccd1 vccd1 _5734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2946_ _2946_/A vssd1 vssd1 vccd1 vccd1 _3144_/A sky130_fd_sc_hd__buf_2
X_5665_ _5694_/CLK _5665_/D vssd1 vssd1 vccd1 vccd1 _5665_/Q sky130_fd_sc_hd__dfxtp_1
X_2877_ _2877_/A vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4988__C _4988_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4616_ _5207_/A vssd1 vssd1 vccd1 vccd1 _4796_/C sky130_fd_sc_hd__buf_2
XFILLER_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4350__A _4350_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5596_ _5641_/CLK _5596_/D vssd1 vssd1 vccd1 vccd1 _5596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5165__B _5178_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3175__A1 _5337_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4478_ _4487_/A _4498_/B _4478_/C vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__or3_1
XFILLER_63_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _3429_/A _3433_/B _4747_/A vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__and3_1
XFILLER_28_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3478__A2 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5181__A _5200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5331__D _5331_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4228__C _4228_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__A1 _5427_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4525__A _4525_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5356__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4898__C _4915_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5506__D _5506_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5312__C1 _5268_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3604__A _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4130__A3 _3994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3874__C1 _3873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3323__B _5552_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output228_A _3318_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5091__A1 _5075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3929__B1 _3918_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ _2800_/A vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__buf_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4051__C1 _4050_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3780_ _3850_/A vssd1 vssd1 vccd1 vccd1 _4283_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3993__B _3993_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2731_ _5751_/Q _2785_/A _2648_/Y _2736_/A vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__o211a_1
XANTENNA__2601__B1 _2600_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5266__A _5266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5450_ _5531_/CLK _5450_/D vssd1 vssd1 vccd1 vccd1 _5450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2662_ _2657_/X _2658_/Y _2613_/X _2661_/Y vssd1 vssd1 vccd1 vccd1 _2748_/B sky130_fd_sc_hd__a31oi_4
XANTENNA__4601__C _4604_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4401_ _5359_/Q _4400_/X _2619_/Y _4379_/X vssd1 vssd1 vccd1 vccd1 _5359_/D sky130_fd_sc_hd__o211a_1
X_5381_ _5765_/CLK _5381_/D vssd1 vssd1 vccd1 vccd1 _5381_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5416__D _5416_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2593_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2904__A1 _2677_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4332_ _4332_/A vssd1 vssd1 vccd1 vccd1 _5329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5303__C1 _5287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4263_ _4263_/A _5308_/A vssd1 vssd1 vccd1 vccd1 _4263_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3514__A _3514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4657__A1 _5478_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3214_ _5196_/C _5344_/Q _3234_/S vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__mux2_8
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2668__B1 _5766_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _5793_/Q _3690_/X _4193_/Y vssd1 vssd1 vccd1 vccd1 _4195_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__4329__B _4333_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3865__C1 _3864_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _5167_/C _5332_/Q _3192_/S vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__mux2_8
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4048__C _4048_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3880__A2 _3879_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3076_ _4542_/B vssd1 vssd1 vccd1 vccd1 _3105_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5082__A1 _5081_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4345__A _4345_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2840__B1 _4411_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4999__B _5005_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3978_ _3978_/A vssd1 vssd1 vccd1 vccd1 _3978_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3396__A1 _5508_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5717_ _5741_/CLK _5717_/D vssd1 vssd1 vccd1 vccd1 _5717_/Q sky130_fd_sc_hd__dfxtp_1
X_2929_ _2929_/A _2929_/B _2929_/C _2929_/D vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__5176__A _5176_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5648_ _5659_/CLK _5648_/D vssd1 vssd1 vccd1 vccd1 _5648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5326__D _5326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5579_ _5694_/CLK _5579_/D vssd1 vssd1 vccd1 vccd1 _5579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4648__A1 _5470_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3424__A _3424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3871__A2 _5002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A ksc_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A1 _5666_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__B2 _5073_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3797__C _3797_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__C1 _4280_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__C1 _4005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input91_A gpio_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4186__B1_N _5477_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3139__A1 _5331_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output178_A _5270_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4887__A1 _4875_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output345_A _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5521__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 cpu_adr_i[15] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4950_ _4950_/A vssd1 vssd1 vccd1 vccd1 _5611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4272__C1 _4271_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5671__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3901_ _4110_/A vssd1 vssd1 vccd1 vccd1 _4079_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2822__B1 _2821_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4881_ _3662_/Y _3678_/X _4847_/X _4191_/Y _4848_/X vssd1 vssd1 vccd1 vccd1 _5581_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3832_ _4082_/A vssd1 vssd1 vccd1 vccd1 _3832_/X sky130_fd_sc_hd__clkbuf_1
X_3763_ _3763_/A vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__buf_2
XANTENNA__3820__A_N _3817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3509__A _3515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5502_ _5538_/CLK _5502_/D vssd1 vssd1 vccd1 vccd1 _5502_/Q sky130_fd_sc_hd__dfxtp_1
X_2714_ _5375_/Q _2621_/X _4431_/B vssd1 vssd1 vccd1 vccd1 _2782_/D sky130_fd_sc_hd__o21ai_2
X_3694_ _4139_/A vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5433_ _5435_/CLK _5433_/D vssd1 vssd1 vccd1 vccd1 _5433_/Q sky130_fd_sc_hd__dfxtp_1
X_2645_ _2645_/A vssd1 vssd1 vccd1 vccd1 _2750_/A sky130_fd_sc_hd__clkbuf_4
Xoutput301 _3523_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[27] sky130_fd_sc_hd__buf_2
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput312 _3481_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4878__A1 _4875_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput323 _3599_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput334 _3635_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5364_ _5800_/CLK _5364_/D vssd1 vssd1 vccd1 vccd1 _5364_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput345 _3566_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2576_ _5261_/A _2616_/A _5261_/D vssd1 vssd1 vccd1 vccd1 _2785_/A sky130_fd_sc_hd__nor3_4
XANTENNA__2889__B1 _2888_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput356 _3002_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput367 _3024_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput378 _2972_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[3] sky130_fd_sc_hd__buf_2
X_4315_ _4439_/C vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__clkbuf_2
Xoutput389 _3130_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5295_ _5295_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5786_/D sky130_fd_sc_hd__nand2_1
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5162__C _5162_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _3824_/A _3857_/A _4244_/X _4245_/X _4835_/A vssd1 vssd1 vccd1 vccd1 _4246_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4082_/X _4083_/X _4177_/C _4257_/D vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__and4bb_1
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3853__A2 _4590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3128_ _4331_/B _5399_/Q _3151_/S vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5055__A1 _5658_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5055__B2 _5034_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3066__A0 _5136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4075__A _4075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3059_ _5133_/C _5318_/Q _4375_/A vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__mux2_8
XFILLER_93_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4803__A _4803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4566__B1 _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4522__B _4526_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5056__D _5056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4869__A1 _4859_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5544__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2696__C _2696_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3154__A _3212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5294__A1 _5785_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__A2 _3954_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5294__B2 _4067_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2993__A _2993_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5694__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5046__A1 _5652_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3601__B _3601_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5046__B2 _5034_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3057__A0 _5703_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__B1 _4425_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4713__A _4713_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4006__C1 _4005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output295_A _3510_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__A2 _5782_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3329__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2887__B _2925_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4190__D1 _3836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3064__A _4617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4100_ _3999_/X _4000_/X _4100_/C _4243_/D vssd1 vssd1 vccd1 vccd1 _4100_/X sky130_fd_sc_hd__and4bb_1
XFILLER_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5080_ _5075_/X _4890_/X _5070_/X _5076_/X _3936_/B vssd1 vssd1 vccd1 vccd1 _5670_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4088__A2 _4080_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__A _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4031_ _3922_/X _3958_/X _3998_/X _4030_/X vssd1 vssd1 vccd1 vccd1 _4031_/X sky130_fd_sc_hd__o211a_1
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3511__B _5650_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3048__A0 _5702_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _5605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4260__A2 _3722_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4623__A _4652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4864_ _4859_/X _4860_/X _4015_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5570_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5417__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3815_ _4489_/A vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__buf_4
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4342__B _4355_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4795_ _5538_/Q _4780_/X _5805_/A _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _5538_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3220__A0 _4366_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3746_ _3869_/A _3746_/B vssd1 vssd1 vccd1 vccd1 _3746_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5157__C _5157_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4217__B_N _3770_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5567__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3677_ _4746_/A _3345_/A _3676_/Y vssd1 vssd1 vccd1 vccd1 _3680_/A sky130_fd_sc_hd__o21ai_2
XFILLER_31_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5416_ _5586_/CLK _5416_/D vssd1 vssd1 vccd1 vccd1 _5416_/Q sky130_fd_sc_hd__dfxtp_1
X_2628_ _2736_/A _2628_/B _2628_/C vssd1 vssd1 vccd1 vccd1 _2628_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__2797__B _2853_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5347_ _5737_/CLK _5347_/D vssd1 vssd1 vccd1 vccd1 _5347_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5604__D _5604_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2559_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__buf_4
XFILLER_62_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput186 _4069_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput197 _4223_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2731__C1 _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3405__C _4729_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5278_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5276__A1 _5771_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5276__B2 _3801_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4229_ _5480_/Q _4489_/A _4228_/X vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3702__A _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4517__B _4526_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4533__A _4533_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4252__B _4252_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3583__S _3597_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input54_A cpu_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5514__D _5514_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4708__A _4708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5019__A1 _5640_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4427__B _4427_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__B2 _5011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output210_A _3949_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output308_A _3472_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A2 _4449_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__B1 _4674_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3600_ _4344_/B _5613_/Q _3600_/S vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__mux2_1
Xinput11 cpu_adr_i[18] vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3202__A0 _5727_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _5433_/D sky130_fd_sc_hd__clkbuf_1
Xinput22 cpu_adr_i[28] vssd1 vssd1 vccd1 vccd1 _2639_/A sky130_fd_sc_hd__clkbuf_2
Xinput33 cpu_adr_i[9] vssd1 vssd1 vccd1 vccd1 _2614_/A sky130_fd_sc_hd__buf_2
Xinput44 cpu_dat_i[18] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3531_ _3531_/A vssd1 vssd1 vccd1 vccd1 _3531_/X sky130_fd_sc_hd__clkbuf_1
Xinput55 cpu_dat_i[28] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
Xinput66 cpu_dat_i[9] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2898__A _4295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput77 gpio_dat_i[12] vssd1 vssd1 vccd1 vccd1 _4001_/C sky130_fd_sc_hd__buf_2
XANTENNA__5274__A _5287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput88 gpio_dat_i[22] vssd1 vssd1 vccd1 vccd1 _4162_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 gpio_dat_i[3] vssd1 vssd1 vccd1 vccd1 _3835_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3462_ _2924_/X _2927_/X _4992_/A vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__o21a_1
X_5201_ _5201_/A vssd1 vssd1 vccd1 vccd1 _5731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3393_ _3393_/A _3397_/B _4722_/A vssd1 vssd1 vccd1 vccd1 _3394_/A sky130_fd_sc_hd__and3_1
XANTENNA__5424__D _5424_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2713__C1 _2637_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5132_ _5156_/A vssd1 vssd1 vccd1 vccd1 _5152_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5258__A1 _5762_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3269__A0 _4390_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5063_ _5068_/A _4664_/A _4252_/C _5204_/A vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__a31o_2
XANTENNA__4618__A _4618_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3522__A _3526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4014_ _3763_/X _3766_/X _3768_/X _4013_/X _3331_/A vssd1 vssd1 vccd1 vccd1 _4014_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4218__C1 _4217_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4233__A2 _4115_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4916_ _4916_/A vssd1 vssd1 vccd1 vccd1 _5599_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3441__A0 _4371_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4353__A _4366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3992__B2 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4847_ _5066_/A vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__buf_4
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4778_ _4778_/A _4778_/B _4778_/C vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__and3_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3744__A1 _3707_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3729_ _4000_/A vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5184__A _5184_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3416__B _3416_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5334__D _5334_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5249__A1 _2696_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4528__A _4528_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4209__C1 _4153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5732__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3432__A0 _4364_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4263__A _4263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2786__A2 _3047_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3983__A1 _3976_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5509__D _5509_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2636__A_N input16/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3607__A _3607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5094__A _5094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output258_A _3417_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4160__A1 _4027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2710__A2 _5261_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4438__A _4438_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5269__A _5289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4215__A2 _4095_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5750_ _5766_/CLK _5750_/D vssd1 vssd1 vccd1 vccd1 _5750_/Q sky130_fd_sc_hd__dfxtp_1
X_2962_ _2876_/X _2882_/X _4548_/A vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4604__C _4604_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4701_ _4701_/A _4707_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__and3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3974__A1 _5464_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5681_ _5697_/CLK _5681_/D vssd1 vssd1 vccd1 vccd1 _5681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5419__D _5419_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2893_ _4098_/A vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__clkbuf_2
X_4632_ _4645_/A vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4901__A _4913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4563_ _4600_/A vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3517__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3514_ _3514_/A vssd1 vssd1 vccd1 vccd1 _3514_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2934__C1 _2779_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4494_ _4514_/A _4498_/B _4494_/C vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__or3_1
XANTENNA__3236__B _4542_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3445_ _3445_/A _3445_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _3446_/A sky130_fd_sc_hd__and3_1
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4151__A1 _4148_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5605__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3376_/A _3380_/B _4709_/C vssd1 vssd1 vccd1 vccd1 _3377_/A sky130_fd_sc_hd__and3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2701__A2 _2683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5115_ _5694_/Q _4913_/B _5060_/X _5114_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _5694_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4348__A _4378_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__C _2794_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5046_ _5652_/Q _5033_/X _5029_/X _5034_/X _5045_/X vssd1 vssd1 vccd1 vccd1 _5652_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5100__B1 _5084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5755__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__B1 _5590_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4206__A2 _3766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5179__A _5179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4083__A _4083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4514__C _4514_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3965__A1 _5779_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3965__B2 _3964_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5329__D _5329_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4811__A _4821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3717__A1 _2728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3427__A _3427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input156_A spi_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4142__B2 _4141_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A cpu_adr_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3653__B1 _4903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4850__C1 _4840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4705__B _4714_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5089__A _5089_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3101__S _3126_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3956__A1 _3956_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4143__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4721__A _4746_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output375_A _2967_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3337__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5628__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5255__C _5264_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2598__D _2684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4118__D1 _4117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2931__A2 _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _4371_/B _5417_/Q _3230_/S vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4133__A1 _3735_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5778__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3161_ _5720_/Q input44/X _3186_/S vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4168__A _4195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5702__D _5702_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3892__B1 _3725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3092_ _3092_/A _3105_/B _4475_/A vssd1 vssd1 vccd1 vccd1 _3093_/A sky130_fd_sc_hd__and3_1
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4436__A2 _2642_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4841__C1 _4840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5802_ _5802_/CLK _5802_/D vssd1 vssd1 vccd1 vccd1 _5802_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3994_ _3994_/A vssd1 vssd1 vccd1 vccd1 _3994_/X sky130_fd_sc_hd__buf_4
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3947__A1 _3813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2945_ _5735_/Q input2/X _3233_/S vssd1 vssd1 vccd1 vccd1 _5210_/C sky130_fd_sc_hd__mux2_2
X_5733_ _5737_/CLK _5733_/D vssd1 vssd1 vccd1 vccd1 _5733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2876_ _3042_/A vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5664_ _5694_/CLK _5664_/D vssd1 vssd1 vccd1 vccd1 _5664_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _5451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5595_ _5641_/CLK _5595_/D vssd1 vssd1 vccd1 vccd1 _5595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4546_ _4546_/A vssd1 vssd1 vccd1 vccd1 _5420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5165__C _5184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4477_ _4558_/B vssd1 vssd1 vccd1 vccd1 _4498_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3428_ _4362_/B _5517_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5181__B _5191_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A cpu_adr_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3359_ _4830_/A vssd1 vssd1 vccd1 vccd1 _3376_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5612__D _5612_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__C1 _3993_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__A _3710_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4541__A _5207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3157__A _3157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2996__A _3042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5312__B1 _5102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5522__D _5522_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3874__B1 _3768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3626__A0 _4360_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4716__A _4716_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3620__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5091__A2 _5089_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3929__A1 _5777_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3929__B2 _3928_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4051__B1 _3975_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4100__B_N _4000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4451__A _4891_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2730_ _2809_/A _2645_/A _5366_/Q vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3993__C _3993_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2601__A1 _5365_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5450__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5266__B _5266_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2661_ _5374_/Q _5376_/Q _2699_/A _2672_/A vssd1 vssd1 vccd1 vccd1 _2661_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4601__D _4614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4400_ _5238_/A vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__buf_4
XFILLER_86_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5380_ _5695_/CLK _5380_/D vssd1 vssd1 vccd1 vccd1 _5380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2592_ input7/X vssd1 vssd1 vccd1 vccd1 _2592_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2904__A2 _5195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4331_ _4344_/A _4331_/B vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__and2_1
XANTENNA__5282__A _5282_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5303__B1 _4193_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4262_ _5798_/Q _3747_/X _4252_/X _4261_/Y vssd1 vssd1 vccd1 vccd1 _5308_/A sky130_fd_sc_hd__o22ai_4
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4657__A2 _4652_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3213_ _5729_/Q input54/X _3223_/S vssd1 vssd1 vccd1 vccd1 _5196_/C sky130_fd_sc_hd__mux2_2
XFILLER_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5432__D _5432_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2668__A1 _2616_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4193_ _5105_/A _3848_/X _4187_/Y _4192_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _4193_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3865__B1 _4835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3192_/S sky130_fd_sc_hd__buf_4
XFILLER_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5067__C1 _3792_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4048__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4626__A _4638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3075_ _3665_/A vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3530__A _3530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5082__A2 _5078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2840__A1 _2839_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3977_ _3977_/A vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4999__C _4999_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5716_ _5741_/CLK _5716_/D vssd1 vssd1 vccd1 vccd1 _5716_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4361__A _4361_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2928_ _2591_/Y _2596_/X _2916_/B _2916_/C vssd1 vssd1 vccd1 vccd1 _2929_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5176__B _5191_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _5659_/CLK _5647_/D vssd1 vssd1 vccd1 vccd1 _5647_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5607__D _5607_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2859_ _5660_/Q vssd1 vssd1 vccd1 vccd1 _2859_/Y sky130_fd_sc_hd__inv_4
XFILLER_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5578_ _5586_/CLK _5578_/D vssd1 vssd1 vccd1 vccd1 _5578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4529_ _4538_/A _4550_/B _4529_/C vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__or3_1
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3705__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5192__A _5192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4648__A2 _4639_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5342__D _5342_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3856__B1 _5087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5323__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__A _4536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3440__A _3440_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A2 _4988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A ksc_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3797__D _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__B1 _5099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5473__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__B1 _4031_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2595__B1 _5749_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input84_A gpio_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5517__D _5517_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4887__A2 _4876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3615__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3772__A_N _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output240_A _3276_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output338_A _3644_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3847__B1 _3846_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4149__C _4149_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5049__C1 _5045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 cpu_adr_i[16] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4446__A _4446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__B1 _3826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3900_ _4240_/A _3900_/B _4240_/C _4240_/D vssd1 vssd1 vccd1 vccd1 _3900_/X sky130_fd_sc_hd__and4_4
XANTENNA__2822__A1 _2817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__A_N _3860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4880_ _4875_/X _4876_/X _4179_/Y _4877_/X vssd1 vssd1 vccd1 vccd1 _5580_/D sky130_fd_sc_hd__a211o_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3831_ _3979_/A vssd1 vssd1 vccd1 vccd1 _3831_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4024__B1 _4023_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_CLK_A clkbuf_1_0_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5277__A _5277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3762_ _3977_/A vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3509__B _5649_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5501_ _5538_/CLK _5501_/D vssd1 vssd1 vccd1 vccd1 _5501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2713_ _2711_/Y _2640_/X _2712_/Y _2637_/A vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__5427__D _5427_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3693_ _5068_/A vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5432_ _5446_/CLK _5432_/D vssd1 vssd1 vccd1 vccd1 _5432_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _5261_/A _5261_/D _2544_/B vssd1 vssd1 vccd1 vccd1 _2645_/A sky130_fd_sc_hd__o21a_1
Xoutput302 _3525_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[28] sky130_fd_sc_hd__buf_2
Xoutput313 _3483_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_86_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4878__A2 _4876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput324 _3602_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[18] sky130_fd_sc_hd__buf_2
X_5363_ _5800_/CLK _5363_/D vssd1 vssd1 vccd1 vccd1 _5363_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput335 _3638_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[28] sky130_fd_sc_hd__buf_2
X_2575_ _5767_/Q vssd1 vssd1 vccd1 vccd1 _2616_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2889__A1 _2886_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput346 _3571_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__3525__A _3525_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput357 _3004_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput368 _3026_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[23] sky130_fd_sc_hd__buf_2
X_4314_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4439_/C sky130_fd_sc_hd__clkbuf_4
Xoutput379 _2978_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[4] sky130_fd_sc_hd__buf_2
X_5294_ _5785_/Q _5289_/X _4058_/X _4067_/Y _5285_/X vssd1 vssd1 vccd1 vccd1 _5785_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5346__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ _3735_/A _4003_/A _5585_/Q vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__o21a_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__B1 _3837_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4176_ _5580_/Q vssd1 vssd1 vccd1 vccd1 _4176_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3127_ _5160_/A _5329_/Q _3162_/S vssd1 vssd1 vccd1 vccd1 _4331_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4356__A _4356_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5055__A2 _5021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5496__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3066__A1 _5319_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3058_ _3144_/A vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4015__B1 _4014_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5187__A _5187_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4566__A1 _5428_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2604__A _2841_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4091__A _4091_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4566__B2 _4564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4522__C _4536_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5337__D _5337_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4869__A2 _4860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5279__C1 _5278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5294__A2 _5289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__A3 _3994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5800__D _5800_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5046__A2 _5033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3601__C _4953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3057__A1 input46/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A1 _2650_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__B1 _4002_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__A _5097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3329__B _5555_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output190_A _3787_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output288_A _3497_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5369__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2887__C _2887_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3345__A _3345_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4190__C1 _4189_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4030_ _3999_/X _4000_/X _4030_/C _4063_/D vssd1 vssd1 vccd1 vccd1 _4030_/X sky130_fd_sc_hd__and4bb_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4176__A _5580_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5710__D _5710_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3048__A1 input35/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4245__B1 _5585_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4904__A _4904_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4932_ _4932_/A _4940_/B _4940_/C vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__and3_1
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _4002_/X _4004_/X _4856_/X _4857_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _5569_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3814_ _4074_/A vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__buf_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4794_ _4794_/A vssd1 vssd1 vccd1 vccd1 _5537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3220__A1 _5415_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3745_ _5769_/Q _3690_/X _3705_/X _3744_/Y vssd1 vssd1 vccd1 vccd1 _3746_/B sky130_fd_sc_hd__o22ai_4
XFILLER_21_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3676_ _3961_/A _3736_/A _5589_/Q vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__o21ai_1
X_5415_ _5531_/CLK _5415_/D vssd1 vssd1 vccd1 vccd1 _5415_/Q sky130_fd_sc_hd__dfxtp_1
X_2627_ _2593_/X _2594_/X _5743_/Q vssd1 vssd1 vccd1 vccd1 _2628_/C sky130_fd_sc_hd__o21ai_2
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2797__C _2797_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4181__C1 _4153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2558_ _5261_/A _5261_/D _2544_/B vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__o21ai_1
X_5346_ _5731_/CLK _5346_/D vssd1 vssd1 vccd1 vccd1 _5346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2731__B1 _2648_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput187 _4090_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput198 _4237_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5277_ _5277_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5772_/D sky130_fd_sc_hd__nand2_1
XANTENNA__5276__A2 _5269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4228_ _4254_/A _4228_/B _4228_/C vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__and3_1
XFILLER_5_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _4240_/A _4159_/B _4159_/C _4214_/D vssd1 vssd1 vccd1 vccd1 _4159_/X sky130_fd_sc_hd__and4_2
XANTENNA__5620__D _5620_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4517__C _4536_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4236__B1 _4226_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4814__A _4821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4252__C _4252_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5511__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2970__A0 _5217_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3165__A _3183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5661__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2722__B1 _2721_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input47_A cpu_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5530__D _5530_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3104__S _3151_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__A2 _5010_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4427__C _4427_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__A _4724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output203_A _4287_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2789__B1 _2916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4242__A3 _3994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__A1 _3281_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4162__C _4162_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3202__A1 input52/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 cpu_adr_i[19] vssd1 vssd1 vccd1 vccd1 _2719_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 cpu_adr_i[29] vssd1 vssd1 vccd1 vccd1 _2697_/A sky130_fd_sc_hd__clkbuf_2
Xinput34 cpu_cyc_i vssd1 vssd1 vccd1 vccd1 _2583_/A sky130_fd_sc_hd__buf_8
Xinput45 cpu_dat_i[19] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_3530_ _3530_/A _5659_/Q vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__and2_1
Xinput56 cpu_dat_i[29] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput67 cpu_sel_i[0] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
Xinput78 gpio_dat_i[13] vssd1 vssd1 vccd1 vccd1 _4013_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2961__A0 _4383_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput89 gpio_dat_i[23] vssd1 vssd1 vccd1 vccd1 _4177_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ _4383_/B _5629_/Q _5033_/A vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5705__D _5705_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3075__A _3665_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5200_/A _5215_/B _5200_/C vssd1 vssd1 vccd1 vccd1 _5201_/A sky130_fd_sc_hd__or3_1
XANTENNA__4163__C1 _4162_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3392_ _4340_/B _5507_/Q _3400_/S vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2713__B1 _2712_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5131_ _5131_/A vssd1 vssd1 vccd1 vccd1 _5702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3803__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5258__A2 _5234_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5062_ _4889_/X _5060_/X _4847_/X _5061_/X _3705_/B vssd1 vssd1 vccd1 vccd1 _5661_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3269__A1 _5528_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3522__B _5655_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4013_ _3860_/X _3861_/X _4013_/C _4278_/D vssd1 vssd1 vccd1 vccd1 _4013_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__5440__D _5440_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4218__B1 _4781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4634__A _4638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4915_ _4915_/A _4915_/B _4915_/C vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__and3_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3441__A1 _5521_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4353__B _4353_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5534__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4846_ _4846_/A vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__buf_2
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4777_ _4777_/A vssd1 vssd1 vccd1 vccd1 _5530_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3744__A2 _4622_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3728_ _4083_/A vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5684__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2952__B1 _4545_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5184__B _5202_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5615__D _5615_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3659_ _3659_/A vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__buf_2
XFILLER_66_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4154__C1 _4153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3416__C _4737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5329_ _5741_/CLK _5329_/D vssd1 vssd1 vccd1 vccd1 _5329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4809__A _4809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5249__A2 _2696_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3713__A _4265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5350__D _5350_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4209__B1 _4208_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4544__A _4678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input101_A gpio_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3432__A1 _5518_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4263__B _5308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3983__A2 _3906_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2999__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5525__D _5525_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4160__A2 _4095_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4719__A _4724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5407__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2710__A3 _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output320_A _3589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output418_A _3241_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3120__A0 _5713_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5557__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4454__A _4454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ _4383_/B _5421_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4604__D _4614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4700_ _4700_/A vssd1 vssd1 vccd1 vccd1 _5498_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3974__A2 _3815_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5680_ _5690_/CLK _5680_/D vssd1 vssd1 vccd1 vccd1 _5680_/Q sky130_fd_sc_hd__dfxtp_1
X_2892_ _2876_/X _2882_/X _3073_/B vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _3756_/X _4667_/C _3853_/Y _3851_/X _4630_/X vssd1 vssd1 vccd1 vccd1 _5457_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4901__B _4913_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3187__A0 _5184_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5285__A _5299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _5427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2934__B1 _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3513_ _3515_/A _5651_/Q vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__and2_1
XANTENNA__5435__D _5435_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4493_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3236__C _4538_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3444_ _4373_/A _5522_/Q _3444_/S vssd1 vssd1 vccd1 vccd1 _4758_/C sky130_fd_sc_hd__mux2_1
XFILLER_63_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3375_ _4329_/A _5502_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _4709_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4151__A2 _4115_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4629__A _5228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3533__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__clkbuf_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5100__A1 _5099_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5045_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3662__A1 _2771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4364__A _4364_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3965__A2 _3915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4829_ _4829_/A vssd1 vssd1 vccd1 vccd1 _5555_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4811__B _5545_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5195__A _5195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3708__A _4128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3717__A2 _3716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5345__D _5345_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4539__A _4539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3443__A _3443_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3350__A0 _4312_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4126__A2_N _5681_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input149_A spi_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3102__A0 _5150_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3653__A1 _3482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4850__B1 _3875_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4705__C _4705_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3956__A2 _3954_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3169__A0 _5176_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3618__A _3618_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output270_A _3352_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output368_A _3026_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4118__C1 _4116_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4251__A1_N _4139_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4133__A2 _4003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__A _4449_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3160_/A vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4168__B _4168_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3892__A1 _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3091_ _4318_/B _5393_/Q _3248_/S vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4841__B1 _3774_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5802_/CLK _5801_/D vssd1 vssd1 vccd1 vccd1 _5801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3993_ _4127_/A _3993_/B _3993_/C _4026_/D vssd1 vssd1 vccd1 vccd1 _3993_/X sky130_fd_sc_hd__and4_2
XFILLER_56_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3947__A2 _3939_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5732_ _5737_/CLK _5732_/D vssd1 vssd1 vccd1 vccd1 _5732_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4912__A _4912_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2944_ _3179_/A vssd1 vssd1 vccd1 vccd1 _3233_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5663_ _5802_/CLK _5663_/D vssd1 vssd1 vccd1 vccd1 _5663_/Q sky130_fd_sc_hd__dfxtp_1
X_2875_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3042_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3528__A _3530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4614_ _4652_/A _5451_/Q _5017_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__and4_1
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5594_ _5641_/CLK _5594_/D vssd1 vssd1 vccd1 vccd1 _5594_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2907__B1 _2906_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4545_ _4674_/A _4550_/B _4545_/C vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__or3_1
XFILLER_85_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3580__A0 _4331_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4476_ _4476_/A vssd1 vssd1 vccd1 vccd1 _5393_/D sky130_fd_sc_hd__clkbuf_1
X_3427_ _3427_/A vssd1 vssd1 vccd1 vccd1 _3427_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4359__A _4385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5722__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3263__A _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5181__C _5181_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3358_ _3358_/A vssd1 vssd1 vccd1 vccd1 _3358_/X sky130_fd_sc_hd__clkbuf_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5085__B1 _5084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4094__A _4127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2607__A _2607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3202__S _3223_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4822__A _4822_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4060__A1 _4027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__A1 _5268_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3874__A1 _3763_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3901__A _4110_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4716__B _4731_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3626__A1 _5620_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3620__B _3620_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5091__A3 _5090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2951__S _3235_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4732__A _4732_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3929__A2 _3915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4051__A1 _3940_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4451__B _4473_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3993__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2601__A2 _2637_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3348__A _3357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5266__C _5266_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2660_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2672_/A sky130_fd_sc_hd__buf_4
XFILLER_86_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2591_ _2569_/X _2704_/A _5364_/Q vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5745__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4330_ _4330_/A vssd1 vssd1 vccd1 vccd1 _5328_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5282__B _5284_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5303__A1 _5793_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _3792_/D _4255_/Y _4260_/Y _4153_/X vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5713__D _5713_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3236_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2668__A2 _2549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4192_ _3824_/X _3857_/X _3826_/X _4191_/Y vssd1 vssd1 vccd1 vccd1 _4192_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3865__A1 _3824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _5717_/Q input41/X _3168_/S vssd1 vssd1 vccd1 vccd1 _5167_/C sky130_fd_sc_hd__mux2_2
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4907__A _4907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5067__B1 _5061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3811__A _4057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3074_ _3074_/A vssd1 vssd1 vccd1 vccd1 _3074_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4626__B _4626_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3530__B _5659_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5082__A3 _5066_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2840__A2 _2762_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4642__A _4651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3976_ _5568_/Q vssd1 vssd1 vccd1 vccd1 _3976_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5715_ _5741_/CLK _5715_/D vssd1 vssd1 vccd1 vccd1 _5715_/Q sky130_fd_sc_hd__dfxtp_1
X_2927_ _2927_/A vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3258__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5646_ _5659_/CLK _5646_/D vssd1 vssd1 vccd1 vccd1 _5646_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5176__C _5176_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2858_ _2845_/X _3664_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3682_/A sky130_fd_sc_hd__o21ai_4
XFILLER_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5577_ _5694_/CLK _5577_/D vssd1 vssd1 vccd1 vccd1 _5577_/Q sky130_fd_sc_hd__dfxtp_1
X_2789_ _2591_/Y _2596_/X _2916_/B vssd1 vssd1 vccd1 vccd1 _2796_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4158__A1_N _3806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3705__B _3705_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4459_ _4459_/A vssd1 vssd1 vccd1 vccd1 _5387_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5623__D _5623_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3856__A1 _3851_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A _4821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3721__A _3755_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__B _4556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__A1 _4628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5618__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3670__B1_N _5694_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__A _4552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4033__A1 _3997_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5230__B1 _2618_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4033__B2 _4032_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5768__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2595__A1 _2593_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input77_A gpio_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2800__A _2800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5533__D _5533_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3847__A1 _5665_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3847__B2 _3847_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4149__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4727__A _4727_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output233_A _3262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3631__A _3631_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5049__B1 _3540_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3935__A1_N _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output400_A _3190_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__A1 _3824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2822__A2 _2642_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3830_ _3978_/A vssd1 vssd1 vccd1 vccd1 _3830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4462__A _4489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4024__B2 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5277__B _5284_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3761_ _4692_/A vssd1 vssd1 vccd1 vccd1 _4743_/A sky130_fd_sc_hd__buf_2
XANTENNA__5708__D _5708_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5500_ _5538_/CLK _5500_/D vssd1 vssd1 vccd1 vccd1 _5500_/Q sky130_fd_sc_hd__dfxtp_1
X_2712_ _2607_/A _2549_/A _5760_/Q vssd1 vssd1 vccd1 vccd1 _2712_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__3783__B1 _3782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3692_ _4138_/A vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5431_ _5435_/CLK _5431_/D vssd1 vssd1 vccd1 vccd1 _5431_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ _5378_/Q _2565_/A _2642_/Y vssd1 vssd1 vccd1 vccd1 _2782_/A sky130_fd_sc_hd__o21ai_4
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3535__A0 _4304_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5293__A _5293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput303 _3527_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__3806__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput314 _5806_/A vssd1 vssd1 vccd1 vccd1 ksc_cyc_o sky130_fd_sc_hd__buf_2
X_5362_ _5800_/CLK _5362_/D vssd1 vssd1 vccd1 vccd1 _5362_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput325 _3607_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2574_ _2574_/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__clkbuf_4
Xoutput336 _3641_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__2889__A2 _4407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput347 _3649_/X vssd1 vssd1 vccd1 vccd1 ksc_sel_o[0] sky130_fd_sc_hd__buf_2
Xoutput358 _3006_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[14] sky130_fd_sc_hd__buf_2
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _5321_/D sky130_fd_sc_hd__clkbuf_1
Xoutput369 _3028_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__5443__D _5443_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5293_ _5293_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5784_/D sky130_fd_sc_hd__nand2_1
X_4244_ _4098_/X _3958_/A _4781_/A _4243_/X vssd1 vssd1 vccd1 vccd1 _4244_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3838__A1 _3827_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4175_ _5476_/Q _4074_/X _4174_/X vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__3541__A _3541_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _5714_/Q input38/X _3126_/S vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__mux2_2
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4799__C1 _4783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3057_ _5703_/Q input46/X _3108_/S vssd1 vssd1 vccd1 vccd1 _5133_/C sky130_fd_sc_hd__mux2_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4372__A _4372_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4015__A1 _4012_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4566__A2 _4563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5618__D _5618_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3959_ _3727_/X _3729_/X _3959_/C _4063_/D vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__and4bb_1
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3774__B1 _3773_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5629_ _5641_/CLK _5629_/D vssd1 vssd1 vccd1 vccd1 _5629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3716__A _4110_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5353__D _5353_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5279__B1 _3867_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4547__A _4595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5440__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input131_A ksc_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3597__S _3597_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A2 _2650_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5590__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A1 _3997_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4006__B2 _4004_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5528__D _5528_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output183_A _4022_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2887__D _2925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4190__B1 _3831_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output350_A _3655_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4457__A _4457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3361__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4245__A1 _3735_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _5604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5288__A _5288_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2705__A _5380_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4862_ _4859_/X _4860_/X _3983_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5568_/D sky130_fd_sc_hd__a211o_1
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3813_ _4059_/A vssd1 vssd1 vccd1 vccd1 _3813_/X sky130_fd_sc_hd__buf_4
XANTENNA__5438__D _5438_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4793_ _4801_/A _5537_/Q _4796_/C vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__and3_1
XFILLER_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4920__A _4938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3744_ _3707_/X _4622_/B _3741_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _3744_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_101_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5313__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3675_ _4098_/A _3957_/A _3961_/A vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__3536__A _3540_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5414_ _5586_/CLK _5414_/D vssd1 vssd1 vccd1 vccd1 _5414_/Q sky130_fd_sc_hd__dfxtp_1
X_2626_ _2695_/C _2695_/D _2836_/A _2695_/B vssd1 vssd1 vccd1 vccd1 _2628_/B sky130_fd_sc_hd__nand4_4
XFILLER_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4181__B1 _4180_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5345_ _5731_/CLK _5345_/D vssd1 vssd1 vccd1 vccd1 _5345_/Q sky130_fd_sc_hd__dfxtp_1
X_2557_ _2581_/A _2583_/A vssd1 vssd1 vccd1 vccd1 _5261_/D sky130_fd_sc_hd__nand2_4
XANTENNA__2731__A1 _5751_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput188 _4106_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[18] sky130_fd_sc_hd__buf_2
XANTENNA__5463__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput199 _4249_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[28] sky130_fd_sc_hd__buf_2
X_5276_ _5771_/Q _5269_/X _3792_/X _3801_/Y _5310_/B vssd1 vssd1 vccd1 vccd1 _5771_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4227_ _4075_/A _4076_/A _4227_/C _4253_/D vssd1 vssd1 vccd1 vccd1 _4228_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__4367__A _4367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _3806_/X _5683_/Q _4157_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _4159_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3109_ _5152_/C _5326_/Q _3132_/S vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__mux2_8
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _5786_/Q _4070_/X _4073_/X _4088_/Y vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__4236__A1 _5796_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4236__B2 _4235_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4814__B _5547_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5198__A _5198_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2615__A _2640_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5348__D _5348_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4252__D _4664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4830__A _4830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3446__A _3446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2970__A1 _5353_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_24_CLK clkbuf_opt_2_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5766_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3165__B _3165_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2722__A1 _5369_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4277__A _5588_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__B _4739_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2789__A1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B1 _3970_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3120__S _3168_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3450__A2 _2899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5336__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output398_A _3178_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3738__B1 _5557_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4740__A _4740_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 cpu_adr_i[1] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
Xinput24 cpu_adr_i[2] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_2
XFILLER_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 cpu_dat_i[0] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_2
Xinput46 cpu_dat_i[1] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 cpu_dat_i[2] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_2
Xinput68 cpu_sel_i[1] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_2
XANTENNA__2961__A1 _5421_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput79 gpio_dat_i[14] vssd1 vssd1 vccd1 vccd1 _4030_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5641_/CLK sky130_fd_sc_hd__clkbuf_16
X_3460_ _3608_/A vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5486__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4163__B1 _4781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3391_ _3391_/A vssd1 vssd1 vccd1 vccd1 _3391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2713__A1 _2711_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5130_/B _5236_/A vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__and3_1
XANTENNA__3910__B1 _3909_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__B _3803_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5112__C1 _5064_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5061_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5721__D _5721_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4012_ _5570_/Q vssd1 vssd1 vccd1 vccd1 _4012_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4915__A _4915_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4218__A1 _4098_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4634__B _4634_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4914_ _4914_/A vssd1 vssd1 vccd1 vccd1 _5598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _4836_/X _4837_/X _3838_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5560_/D sky130_fd_sc_hd__a211o_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4776_ _4913_/A _4776_/B _4776_/C vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__or3_1
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3727_ _3999_/A vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2952__A1 _2876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5184__C _5184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3658_ _2726_/A _3666_/A _2845_/X vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__a21oi_4
XFILLER_88_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4154__B1 _4152_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2609_ input5/X vssd1 vssd1 vccd1 vccd1 _2610_/A sky130_fd_sc_hd__inv_2
XFILLER_66_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3589_ _3589_/A vssd1 vssd1 vccd1 vccd1 _3589_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5328_ _5741_/CLK _5328_/D vssd1 vssd1 vccd1 vccd1 _5328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5103__C1 _4159_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5631__D _5631_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5259_ _2639_/Y _5227_/X _2641_/Y _4848_/A _4429_/X vssd1 vssd1 vccd1 vccd1 _5763_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4825__A _4828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4209__A1 _3792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5359__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3968__B1 _3967_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4560__A _4711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2999__B _5431_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4719__B _4739_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5541__D _5541_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3115__S _3162_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3120__A1 input37/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output313_A _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4735__A _4971_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5482_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4454__B _4475_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2960_ _3252_/S vssd1 vssd1 vccd1 vccd1 _3240_/S sky130_fd_sc_hd__buf_2
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4173__C _4173_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _3196_/A vssd1 vssd1 vccd1 vccd1 _3073_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4470__A _4470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4630_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__buf_4
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4901__C _4901_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3187__A1 _5339_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4561_ _4561_/A _4681_/B _4569_/A vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__and3_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5716__D _5716_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2934__A1 _4439_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3512_ _3512_/A vssd1 vssd1 vccd1 vccd1 _3512_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ _4492_/A vssd1 vssd1 vccd1 vccd1 _5399_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4136__B1 _4127_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3443_ _3443_/A vssd1 vssd1 vccd1 vccd1 _3443_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3814__A _4074_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A vssd1 vssd1 vccd1 vccd1 _3374_/X sky130_fd_sc_hd__clkbuf_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3895__C1 _3743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5099_/X _5094_/A _5066_/A _5102_/X _3674_/A vssd1 vssd1 vccd1 vccd1 _5693_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__D _5451_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5044_ _5044_/A vssd1 vssd1 vccd1 vccd1 _5651_/D sky130_fd_sc_hd__clkbuf_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5100__A2 _5094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5501__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4645__A _4645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3662__A2 _3998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2870__B1 _5268_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4364__B _4381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5651__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4828_ _4828_/A _5555_/Q _4988_/C vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__and3_1
XANTENNA__4811__C _4817_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4759_ _4759_/A vssd1 vssd1 vccd1 vccd1 _5522_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5626__D _5626_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3724__A _3998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2689__B1 _2688_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3350__A1 _5495_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5361__D _5361_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3102__A1 _5325_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__A _4555_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3653__A2 _2927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4850__A1 _4836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5260__D1 _4377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3956__A3 _3714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4290__A _4378_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3169__A1 _5336_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5536__D _5536_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4118__B1 _3979_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output263_A _3434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3634__A _3646_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5524__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3892__A2 _3723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3090_ _5145_/A _5323_/Q _3102_/S vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4465__A _4465_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4841__A1 _4836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5674__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5800_ _5800_/CLK _5800_/D vssd1 vssd1 vccd1 vccd1 _5800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3989_/X _5673_/Q _3990_/Y _3991_/X vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5731_ _5731_/CLK _5731_/D vssd1 vssd1 vccd1 vccd1 _5731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2943_ _3047_/A vssd1 vssd1 vccd1 vccd1 _3179_/A sky130_fd_sc_hd__buf_2
XANTENNA__3801__C1 _3743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5662_ _5692_/CLK _5662_/D vssd1 vssd1 vccd1 vccd1 _5662_/Q sky130_fd_sc_hd__dfxtp_1
X_2874_ _5452_/Q vssd1 vssd1 vccd1 vccd1 _3029_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3528__B _5658_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4613_ _5450_/Q _4573_/D _3062_/A _4590_/A _4598_/X vssd1 vssd1 vccd1 vccd1 _5450_/D
+ sky130_fd_sc_hd__a221o_1
X_5593_ _5641_/CLK _5593_/D vssd1 vssd1 vccd1 vccd1 _5593_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5446__D _5446_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2907__A1 _2826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4544_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3580__A1 _5607_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4475_ _4475_/A _4475_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__and3_1
XANTENNA__3544__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3426_ _3429_/A _3433_/B _4744_/C vssd1 vssd1 vccd1 vccd1 _3427_/A sky130_fd_sc_hd__and3_1
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3357_ _3357_/A _3361_/B _4697_/A vssd1 vssd1 vccd1 vccd1 _3358_/A sky130_fd_sc_hd__and3_1
XFILLER_24_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4078__C _4078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3288_ _3292_/A _5536_/Q vssd1 vssd1 vccd1 vccd1 _3289_/A sky130_fd_sc_hd__and2_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5085__A1 _5081_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5043_/A _5643_/Q _5039_/C _5043_/D vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__and4_1
XANTENNA__3096__A0 _5148_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4375__A _4375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4094__B _4094_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4060__A2 _3919_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3719__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2623__A _2647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5356__D _5356_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5547__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input161_A spi_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5312__A2 _5096_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3874__A2 _3766_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5697__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input22_A cpu_adr_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4716__C _4716_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3620__C _4963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5233__D1 _4377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4051__A2 _4046_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4451__C _4451_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3348__B _3361_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output380_A _2982_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3853__B1_N _5457_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2590_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__buf_4
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4147_/X _3722_/X _3758_/A _4259_/Y vssd1 vssd1 vccd1 vccd1 _4260_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5303__A2 _5114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3211_ _3211_/A vssd1 vssd1 vccd1 vccd1 _3211_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4188_/Y _3828_/X _4190_/Y vssd1 vssd1 vccd1 vccd1 _4191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3865__A2 _3857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3142_ _3142_/A vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4907__B _4915_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5067__A1 _4889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3078__A0 _5706_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4195__A _4195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3073_ _3092_/A _3073_/B _4469_/C vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__and3_1
XFILLER_3_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2708__A _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2825__B1 _4431_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4923__A _5025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4642__B _4642_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3975_ _4005_/A vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5714_ _5766_/CLK _5714_/D vssd1 vssd1 vccd1 vccd1 _5714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3250__A0 _5701_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2926_ _4295_/D vssd1 vssd1 vccd1 vccd1 _2927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4001__A_N _3999_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5645_ _5659_/CLK _5645_/D vssd1 vssd1 vccd1 vccd1 _5645_/Q sky130_fd_sc_hd__dfxtp_1
X_2857_ _2560_/Y _2949_/A _5802_/Q vssd1 vssd1 vccd1 vccd1 _3669_/B sky130_fd_sc_hd__a21oi_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5576_ _5586_/CLK _5576_/D vssd1 vssd1 vccd1 vccd1 _5576_/Q sky130_fd_sc_hd__dfxtp_1
X_2788_ _2788_/A _2788_/B vssd1 vssd1 vccd1 vccd1 _2853_/C sky130_fd_sc_hd__nor2_4
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _5413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _4458_/A _4475_/B _4542_/A vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__and3_1
XANTENNA__3705__C _5090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3409_ _3412_/A _3416_/B _4731_/A vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__and3_1
XFILLER_28_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _5353_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3856__A2 _3853_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__B _5549_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3213__S _3223_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4536__C _4536_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__A2 _3857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4833__A _5087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__B _4556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5230__A1 _2614_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4033__A2 _3890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3241__B1 _4445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2595__A2 _2594_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3184__A _3184_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3847__A2 _4986_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5049__A1 _5654_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5049__B2 _5034_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output226_A _3313_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__A2_N _5669_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__B1 _5381_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4272__A2 _3825_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4743__A _4743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_1_CLK clkbuf_1_1_1_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_CLK/X sky130_fd_sc_hd__clkbuf_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3359__A _4830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5712__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _4115_/A vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _2711_/A vssd1 vssd1 vccd1 vccd1 _2711_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3783__A1 _5454_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3691_ _5694_/Q _4968_/A _2870_/Y vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__o21a_1
XFILLER_88_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5430_ _5435_/CLK _5430_/D vssd1 vssd1 vccd1 vccd1 _5430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _2639_/Y _2640_/X _2641_/Y _2574_/A vssd1 vssd1 vccd1 vccd1 _2642_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_86_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3535__A1 _5595_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5293__B _5297_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput304 _3464_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[2] sky130_fd_sc_hd__buf_2
X_5361_ _5800_/CLK _5361_/D vssd1 vssd1 vccd1 vccd1 _5361_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4193__D1 _3866_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput315 _3537_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[0] sky130_fd_sc_hd__buf_2
X_2573_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__clkbuf_4
Xoutput326 _3541_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__3094__A _4617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5724__D _5724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput337 _3545_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_86_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4312_ _4322_/A _4312_/B vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__and2_1
XANTENNA__2743__C1 _2637_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput348 _3651_/X vssd1 vssd1 vccd1 vccd1 ksc_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_86_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput359 _3009_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[15] sky130_fd_sc_hd__buf_2
X_5292_ _5783_/Q _5289_/X _4026_/X _4034_/Y _5285_/X vssd1 vssd1 vccd1 vccd1 _5783_/D
+ sky130_fd_sc_hd__o221a_1
X_4243_ _3769_/X _3770_/X _4243_/C _4243_/D vssd1 vssd1 vccd1 vccd1 _4243_/X sky130_fd_sc_hd__and4bb_1
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4918__A _4968_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3838__A2 _3828_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4254_/A _4228_/B _4174_/C vssd1 vssd1 vccd1 vccd1 _4174_/X sky130_fd_sc_hd__and3_1
XFILLER_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4799__B1 _4798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3056_ _3179_/A vssd1 vssd1 vccd1 vccd1 _3108_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3471__A0 _4390_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5392__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4015__A2 _4743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3223__A0 _5731_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4420__C1 _4299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _3958_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3774__A1 _3759_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2909_ _2909_/A _2909_/B _2909_/C _2929_/B vssd1 vssd1 vccd1 vccd1 _2910_/C sky130_fd_sc_hd__nand4_1
X_3889_ _3889_/A1 _4528_/A _3714_/X _3888_/Y vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__a31oi_4
XANTENNA__2901__A _2935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5628_ _5692_/CLK _5628_/D vssd1 vssd1 vccd1 vccd1 _5628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5559_ _5802_/CLK _5559_/D vssd1 vssd1 vccd1 vccd1 _5559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5634__D _5634_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3208__S _3219_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5279__A1 _5773_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4828__A _4828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input124_A ksc_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5735__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4563__A _4600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3462__B1 _4992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A2 _3890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3179__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__A0 _5196_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5544__D _5544_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4190__A1 _3829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_0_CLK CLK vssd1 vssd1 vccd1 vccd1 clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_83_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4738__A _4738_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output343_A _3559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4142__A1_N _4139_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3361__B _3361_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4245__A2 _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3453__A0 _4301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4473__A _4487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4930_ _4938_/A _4938_/B _4930_/C vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__or3_1
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4650__C1 _4645_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5288__B _5297_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4861_ _5268_/A vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5719__D _5719_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3812_ _4240_/A _3812_/B _4240_/C _4240_/D vssd1 vssd1 vccd1 vccd1 _3812_/X sky130_fd_sc_hd__and4_4
X_4792_ _5536_/Q _4780_/X _5805_/A _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _5536_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3902__B_N _3818_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3743_ _4070_/A vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4920__B _4938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3817__A _4075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3674_ _3674_/A _3682_/A _3790_/A vssd1 vssd1 vccd1 vccd1 _3681_/C sky130_fd_sc_hd__nand3_1
XANTENNA__3536__B _3547_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5413_ _5531_/CLK _5413_/D vssd1 vssd1 vccd1 vccd1 _5413_/Q sky130_fd_sc_hd__dfxtp_1
X_2625_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2695_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5454__D _5454_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3809__A2_N _5664_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4181__A1 _4042_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5344_ _5731_/CLK _5344_/D vssd1 vssd1 vccd1 vccd1 _5344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5608__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2556_ _5768_/Q vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput178 _5270_/B vssd1 vssd1 vccd1 vccd1 cpu_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__2731__A2 _2785_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput189 _4123_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[19] sky130_fd_sc_hd__buf_2
X_5275_ _5275_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5770_/D sky130_fd_sc_hd__nand2_1
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3552__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4226_ _4252_/A _4226_/B _4252_/C _4664_/A vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__and4_4
XFILLER_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5758__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4157_ _4157_/A vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3108_ _5711_/Q input66/X _3108_/S vssd1 vssd1 vccd1 vccd1 _5152_/C sky130_fd_sc_hd__mux2_2
XFILLER_99_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _4042_/X _4080_/Y _4087_/Y _3946_/X vssd1 vssd1 vccd1 vccd1 _4088_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__4236__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3039_ _3039_/A vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3444__A0 _4373_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4383__A _4396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4814__C _4817_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3907__A_N _3832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5198__B _5202_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3995__A1 _3794_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5629__D _5629_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4830__B _4830_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3727__A _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5364__D _5364_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3165__C _4508_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2722__A2 _2565_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4558__A _4674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4880__C1 _4877_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__A0 _4366_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4293__A _4293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2806__A _2806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4724__C _4724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2789__A2 _2596_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3986__A1 _5780_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B2 _3985_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5539__D _5539_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3738__A1 _4830_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output293_A _3462_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3637__A _3646_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput14 cpu_adr_i[20] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 cpu_adr_i[30] vssd1 vssd1 vccd1 vccd1 _5261_/C sky130_fd_sc_hd__buf_4
Xinput36 cpu_dat_i[10] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2541__A input3/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput47 cpu_dat_i[20] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput58 cpu_dat_i[30] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 cpu_sel_i[2] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4163__A1 _4098_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3390_ _3393_/A _3397_/B _4719_/C vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__and3_1
XANTENNA__2713__A2 _2640_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3910__A1 _3905_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4468__A _4678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5060_ _5094_/A vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5112__B1 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _5674_/Q _5002_/A _3846_/X _5086_/B2 vssd1 vssd1 vccd1 vccd1 _4011_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4871__C1 _4861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4915__B _4915_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4218__A2 _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5299__A _5299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4913_ _4913_/A _4913_/B _4913_/C vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__or3_1
XANTENNA__5449__D _5449_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4931__A _4931_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4844_ _3798_/X _3799_/X _4832_/X _4833_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _5559_/D
+ sky130_fd_sc_hd__o221a_1
X_4775_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__buf_4
XANTENNA__3547__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3726_ _4082_/A vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5430__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2952__A2 _2882_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3657_ _3711_/A _2854_/X _2845_/X vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4154__A1 _4042_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2608_ _2607_/X _2549_/X _5747_/Q vssd1 vssd1 vccd1 vccd1 _2611_/B sky130_fd_sc_hd__o21bai_1
X_3588_ _3594_/A _3601_/B _4940_/A vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__and3_1
XANTENNA__5580__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2539_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2691_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4378__A _4378_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5327_ _5741_/CLK _5327_/D vssd1 vssd1 vccd1 vccd1 _5327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3282__A _3282_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5103__B1 _5102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5762_/Q _5234_/A _2819_/Y _5228_/X _4377_/X vssd1 vssd1 vccd1 vccd1 _5762_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4209_ _3792_/D _4203_/Y _4208_/Y _4153_/X vssd1 vssd1 vccd1 vccd1 _4209_/Y sky130_fd_sc_hd__o211ai_2
X_5189_ _5189_/A _5202_/B _5208_/C vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__and3_1
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4862__C1 _4861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4825__B _5553_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4209__A2 _4203_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2626__A _2695_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5002__A _5002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3968__B2 _3934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5359__D _5359_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2928__C1 _2916_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input52_A cpu_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4288__A input1/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4719__C _4719_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3656__B1 _5268_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4853__C1 _4843_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3408__A0 _4349_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output306_A _3531_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3131__S _3168_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4454__C _4542_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4173__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2970__S _3229_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4751__A _4751_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2890_ _3665_/A vssd1 vssd1 vccd1 vccd1 _3196_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5453__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5030__C1 _5023_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3367__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4253__B_N _4076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3511_ _3515_/A _5650_/Q vssd1 vssd1 vccd1 vccd1 _3512_/A sky130_fd_sc_hd__and2_1
XANTENNA__2934__A2 _4439_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4491_ _4491_/A _4500_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__and3_1
XFILLER_85_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4136__A1 _5789_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3442_ _3445_/A _3445_/B _4756_/A vssd1 vssd1 vccd1 vccd1 _3443_/A sky130_fd_sc_hd__and3_1
XANTENNA__4136__B2 _4135_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3373_ _3376_/A _3380_/B _4707_/A vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__and3_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5732__D _5732_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__B1 _3894_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5112_ _5692_/Q _4988_/A _3750_/X _5112_/B2 _5064_/A vssd1 vssd1 vccd1 vccd1 _5692_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5043_ _5043_/A _5651_/Q _5056_/C _5043_/D vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__and4_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4926__A _4938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5100__A3 _5087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3830__A _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__C1 _4843_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2870__A1 _2861_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4072__B1 _4071_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4827_ _5554_/Q _4803_/A _3339_/A _4804_/A _4823_/X vssd1 vssd1 vccd1 vccd1 _5554_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3277__A _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4758_ _4771_/A _4763_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__or3_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3709_ _3709_/A vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__clkbuf_2
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _5494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5642__D _5642_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2689__A1 _2682_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5088__C1 _4026_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5326__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4836__A _5081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3740__A _4005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4850__A2 _4837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5476__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5260__C1 _5228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5012__C1 _4823_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3915__A _4091_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4118__A1 _3977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3634__B _3637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5552__D _5552_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output256_A _3410_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3126__S _3126_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__B1 _3876_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5079__C1 _3918_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2965__S _3251_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4746__A _4746_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3629__A0 _4362_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output423_A _2892_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4841__A2 _4837_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _4141_/A vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__buf_2
XANTENNA__5251__C1 _5238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4481__A _4481_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5730_ _5731_/CLK _5730_/D vssd1 vssd1 vccd1 vccd1 _5730_/Q sky130_fd_sc_hd__dfxtp_1
X_2942_ _2924_/X _2927_/X _3547_/B vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3801__B1 _3800_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5661_ _5802_/CLK _5661_/D vssd1 vssd1 vccd1 vccd1 _5661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2873_ _2776_/Y _3790_/A _3682_/A _3683_/A _5268_/C vssd1 vssd1 vccd1 vccd1 _5270_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__5727__D _5727_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3097__A _3163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4612_ _4612_/A vssd1 vssd1 vccd1 vccd1 _5449_/D sky130_fd_sc_hd__clkbuf_1
X_5592_ _5635_/CLK _5592_/D vssd1 vssd1 vccd1 vccd1 _5592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2907__A2 _2717_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4543_ _4543_/A vssd1 vssd1 vccd1 vccd1 _5419_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3825__A _3857_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _5392_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3544__B _3547_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5349__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3425_ _4360_/A _5516_/Q _3432_/S vssd1 vssd1 vccd1 vccd1 _4744_/C sky130_fd_sc_hd__mux2_1
XFILLER_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5462__D _5462_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3868__B1 _3867_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3356_ _4318_/B _5497_/Q _3364_/S vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4149__B_N _4083_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4078__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3287_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3287_/X sky130_fd_sc_hd__clkbuf_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__A _5058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5499__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5085__A2 _5078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3096__A1 _5324_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2843__A1 _5696_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4094__C _4159_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4045__B1 _4044_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4391__A _4391_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5637__D _5637_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3735__A _3735_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5372__D _5372_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5312__A3 _5114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4269__C _4269_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input154_A spi_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3470__A _4295_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4284__B1 _4283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input15_A cpu_adr_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5233__C1 _5228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5547__D _5547_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3348__C _4688_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output373_A _3037_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5303__A3 _5069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3210_ _3210_/A _3221_/B _4526_/A vssd1 vssd1 vccd1 vccd1 _3211_/A sky130_fd_sc_hd__and3_1
XFILLER_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5641__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4190_ _3829_/X _3830_/X _3831_/X _4189_/X _3836_/X vssd1 vssd1 vccd1 vccd1 _4190_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3141_ _3152_/A _3165_/B _4496_/A vssd1 vssd1 vccd1 vccd1 _3142_/A sky130_fd_sc_hd__and3_1
XANTENNA__4476__A _4476_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3380__A _3393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4907__C _4915_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5067__A2 _5060_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _4310_/A _5390_/Q _3230_/S vssd1 vssd1 vccd1 vccd1 _4469_/C sky130_fd_sc_hd__mux2_1
XFILLER_97_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3078__A1 input61/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4195__B _4195_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5791__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2825__A1 _2823_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2825__B2 _4431_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2695__A_N input14/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2724__A _2724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3974_ _5464_/Q _3815_/X _3973_/X vssd1 vssd1 vccd1 vccd1 _3974_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_91_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5713_ _5765_/CLK _5713_/D vssd1 vssd1 vccd1 vccd1 _5713_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3250__A1 input70/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2925_ _2925_/A _2925_/B _2925_/C vssd1 vssd1 vccd1 vccd1 _4295_/D sky130_fd_sc_hd__and3_4
XANTENNA__5457__D _5457_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5644_ _5659_/CLK _5644_/D vssd1 vssd1 vccd1 vccd1 _5644_/Q sky130_fd_sc_hd__dfxtp_1
X_2856_ _2561_/Y _2949_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _3664_/A sky130_fd_sc_hd__a21oi_2
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5575_ _5694_/CLK _5575_/D vssd1 vssd1 vccd1 vccd1 _5575_/Q sky130_fd_sc_hd__dfxtp_1
X_2787_ _2787_/A _2787_/B _2787_/C _2935_/B vssd1 vssd1 vccd1 vccd1 _2788_/B sky130_fd_sc_hd__nand4_2
XANTENNA__3555__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4526_ _4526_/A _4526_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__and3_1
XFILLER_85_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4457_ _4457_/A vssd1 vssd1 vccd1 vccd1 _5386_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3705__D _3792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3408_ _4349_/B _5511_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4388_ _4396_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__and2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A cpu_adr_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3339_ _3339_/A _4761_/A _4683_/C vssd1 vssd1 vccd1 vccd1 _3340_/A sky130_fd_sc_hd__and3_1
XFILLER_24_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__A _4386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3290__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__C _4817_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2634__A _2684_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5010__A _5056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4552__C _4569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5230__A2 _5227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3241__A1 _2973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5367__D _5367_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5514__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3465__A _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5664__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2752__B1 _2751_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2809__A _2809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4296__A _4385_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3404__S _3432_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5049__A2 _5033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__A1 _2806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output219_A _3300_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4009__B1 _3993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2544__A _2544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4060__B1_N _5469_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2710_ _5261_/B _5261_/C _2708_/X _2709_/Y _2606_/X vssd1 vssd1 vccd1 vccd1 _4439_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3783__A2 _4444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3690_ _4091_/A vssd1 vssd1 vccd1 vccd1 _3690_/X sky130_fd_sc_hd__buf_4
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2641_ _2616_/X _2617_/X _5763_/Q vssd1 vssd1 vccd1 vccd1 _2641_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__4193__C1 _4192_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput305 _3529_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[30] sky130_fd_sc_hd__buf_2
X_2572_ _5363_/Q vssd1 vssd1 vccd1 vccd1 _2572_/Y sky130_fd_sc_hd__inv_2
X_5360_ _5800_/CLK _5360_/D vssd1 vssd1 vccd1 vccd1 _5360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput316 _3575_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput327 _3611_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__2743__B1 _2742_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput338 _3644_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[30] sky130_fd_sc_hd__buf_2
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _5320_/D sky130_fd_sc_hd__clkbuf_1
Xoutput349 _3653_/X vssd1 vssd1 vccd1 vccd1 ksc_sel_o[2] sky130_fd_sc_hd__buf_2
X_5291_ _5291_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5782_/D sky130_fd_sc_hd__nand2_1
XFILLER_64_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4242_ _4242_/A1 _4449_/A _3994_/A _4241_/Y vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__a31oi_4
XFILLER_25_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _4075_/X _4076_/X _4173_/C _4201_/D vssd1 vssd1 vccd1 vccd1 _4174_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__5740__D _5740_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2719__A _2719_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3124_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4248__B1 _4240_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _3055_/A vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4799__A1 _5540_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4799__B2 _4782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4934__A _4938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3981__B_N _3833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3471__A1 _5632_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5537__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3223__A1 input56/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4028__B1_N _5467_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4420__B1 _2721_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2908_ _2908_/A _2908_/B _2908_/C _2908_/D vssd1 vssd1 vccd1 vccd1 _2910_/B sky130_fd_sc_hd__nand4_2
XANTENNA__3774__A2 _4743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3888_ _3794_/X _3716_/X _5459_/Q vssd1 vssd1 vccd1 vccd1 _3888_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__5687__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2982__B1 _4556_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5627_ _5697_/CLK _5627_/D vssd1 vssd1 vccd1 vccd1 _5627_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2901__B _2935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2839_ _2809_/X _2750_/X _5361_/Q vssd1 vssd1 vccd1 vccd1 _2839_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3285__A _3285_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5558_ _5589_/CLK _5558_/D vssd1 vssd1 vccd1 vccd1 _5558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4509_ _4509_/A vssd1 vssd1 vccd1 vccd1 _5405_/D sky130_fd_sc_hd__clkbuf_1
X_5489_ _5531_/CLK _5489_/D vssd1 vssd1 vccd1 vccd1 _5489_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5279__A2 _5114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4828__B _5555_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5650__D _5650_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3224__S _3234_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5005__A _5128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4239__B1 _4238_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A ksc_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3462__A1 _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3214__A1 _5344_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input82_A gpio_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3195__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__B1 _2561_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4190__A2 _3830_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3923__A _4099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2539__A _2621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output336_A _3641_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5560__D _5560_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3150__A0 _5169_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3361__C _4699_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4754__A _4771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4473__B _4473_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3453__A1 _5490_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4650__B1 _4112_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4860_ _5089_/A vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3811_ _4057_/A vssd1 vssd1 vccd1 vccd1 _4240_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4791_ _4791_/A vssd1 vssd1 vccd1 vccd1 _5535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3742_ _3742_/A vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__buf_2
XANTENNA__4920__C _4920_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5735__D _5735_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3673_ _4139_/A _3549_/A _3672_/Y vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__4166__C1 _3840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5412_ _5586_/CLK _5412_/D vssd1 vssd1 vccd1 vccd1 _5412_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3536__C _4907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2624_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2695_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2716__B1 _5753_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4181__A2 _4175_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5343_ _5731_/CLK _5343_/D vssd1 vssd1 vccd1 vccd1 _5343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4929__A _4929_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2555_ _2809_/A vssd1 vssd1 vccd1 vccd1 _2675_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3833__A _4083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput179 _3746_/Y vssd1 vssd1 vccd1 vccd1 cpu_dat_o[0] sky130_fd_sc_hd__buf_2
X_5274_ _5287_/A vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3552__B _3565_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4225_ _4139_/X _5688_/Q _4224_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_29_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5470__D _5470_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4156_ _4195_/A _5300_/A vssd1 vssd1 vccd1 vccd1 _4156_/Y sky130_fd_sc_hd__nor2_4
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3107_ _3196_/A vssd1 vssd1 vccd1 vccd1 _3134_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4664__A _4664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4087_ _3940_/X _4046_/X _3975_/X _4086_/Y vssd1 vssd1 vccd1 vccd1 _4087_/Y sky130_fd_sc_hd__o211ai_1
X_3038_ _3038_/A _5449_/Q vssd1 vssd1 vccd1 vccd1 _3039_/A sky130_fd_sc_hd__and2_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3444__A1 _5522_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4383__B _4383_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3995__A2 _3919_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5198__C _5208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4830__C _4988_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2955__A0 _5736_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5645__D _5645_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2631__B _2909_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3219__S _3219_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4839__A _5097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3743__A _4070_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_CLK clkbuf_1_0_1_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4558__B _4558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5380__D _5380_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5702__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3132__A0 _5162_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4880__B1 _4179_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4574__A _4574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__A1 _5519_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__A2 _3804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3199__A0 _4357_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3918__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3738__A2 _3737_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3637__B _3637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput15 cpu_adr_i[21] vssd1 vssd1 vccd1 vccd1 _2663_/C sky130_fd_sc_hd__buf_2
Xinput26 cpu_adr_i[31] vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5555__D _5555_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output286_A _3492_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput37 cpu_dat_i[11] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 cpu_dat_i[21] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput59 cpu_dat_i[31] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4163__A2 _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4749__A _4749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3910__A2 _3906_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5382__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5112__A1 _5692_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5112__B2 _5112_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4010_ _4036_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4010_/Y sky130_fd_sc_hd__nor2_8
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4871__B1 _4119_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4484__A _4484_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4915__C _4915_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _4912_/A vssd1 vssd1 vccd1 vccd1 _5597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4843_ _5235_/A vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3828__A _4692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4774_ _4774_/A vssd1 vssd1 vccd1 vccd1 _5529_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3547__B _3547_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3725_ _4781_/A vssd1 vssd1 vccd1 vccd1 _3725_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5465__D _5465_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3656_ _2560_/Y _2949_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__a21o_2
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2607_ _2607_/A vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4154__A2 _4146_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3587_ _4335_/B _5609_/Q _3600_/S vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5725__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3563__A _3563_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5326_ _5695_/CLK _5326_/D vssd1 vssd1 vccd1 vccd1 _5326_/Q sky130_fd_sc_hd__dfxtp_1
X_2538_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2570__D1 _2569_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5103__A1 _5099_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5257_ _2783_/X _2671_/Y _4565_/X _4400_/X vssd1 vssd1 vccd1 vccd1 _5761_/D sky130_fd_sc_hd__a211o_1
X_4208_ _4147_/X _3722_/X _3758_/A _4207_/Y vssd1 vssd1 vccd1 vccd1 _4208_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5188_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5208_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__4862__B1 _3983_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4394__A _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4139_ _4139_/A vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__buf_4
XFILLER_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4825__C _4988_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2626__B _2695_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2928__B1 _2916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5375__D _5375_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4569__A _4569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3353__A0 _4316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input45_A cpu_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3656__A1 _2560_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4853__B1 _4832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3408__A1 _5511_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__B _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output201_A _3803_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4751__B _4756_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5030__B1 _5029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5748__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3510_ _3510_/A vssd1 vssd1 vccd1 vccd1 _3510_/X sky130_fd_sc_hd__clkbuf_1
X_4490_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4512_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _4371_/B _5521_/Q _3441_/S vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4136__A2 _4091_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4479__A _4479_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3372_ _4327_/B _5501_/Q _3400_/S vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__A1 _3887_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _5111_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5691_/D sky130_fd_sc_hd__nor2_1
XFILLER_83_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5056_/C sky130_fd_sc_hd__clkbuf_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4926__B _4938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__B1 _4832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2727__A _3849_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2870__A2 _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4942__A _5270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4072__B2 _3934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3558__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4826_ _4826_/A vssd1 vssd1 vccd1 vccd1 _5553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4078__B_N _4076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4757_ _4757_/A vssd1 vssd1 vccd1 vccd1 _5521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3583__A0 _4333_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3708_ _4128_/A vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4688_ _4699_/A _4688_/B _4688_/C vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__or3_1
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3639_ _4368_/A _5624_/Q _3645_/S vssd1 vssd1 vccd1 vccd1 _4980_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4389__A _4389_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3293__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2689__A2 _2565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5309_ _5799_/Q _5114_/A _5069_/X _4273_/Y _5287_/A vssd1 vssd1 vccd1 vccd1 _5799_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5088__B1 _5084_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2637__A _2637_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5013__A _5033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4599__C1 _4598_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5260__B1 _2698_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5012__B1 _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4118__A2 _3978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4299__A _4299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3634__C _4976_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3877__A1 _3871_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output249_A _3388_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5079__B1 _5061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__A _4138_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3629__A1 _5621_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output416_A _3106_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2837__C1 _2696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2547__A _2607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5420__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2981__S _3240_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4762__A _4762_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3990_ _3990_/A vssd1 vssd1 vccd1 vccd1 _3990_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5251__B1 _4891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2941_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3547_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4481__B _4500_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3801__A1 _3707_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3378__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5570__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5660_ _5694_/CLK _5660_/D vssd1 vssd1 vccd1 vccd1 _5660_/Q sky130_fd_sc_hd__dfxtp_4
X_2872_ _5261_/B _5261_/D _2544_/A vssd1 vssd1 vccd1 vccd1 _5268_/C sky130_fd_sc_hd__o21a_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4611_ _4611_/A _5449_/Q _5017_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4612_/A sky130_fd_sc_hd__and4_1
XFILLER_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5591_ _5641_/CLK _5591_/D vssd1 vssd1 vccd1 vccd1 _5591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4542_ _4542_/A _4542_/B _5266_/B vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__and3_1
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4473_ _4487_/A _4473_/B _4473_/C vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__or3_1
XANTENNA__5743__D _5743_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3424_ _3424_/A vssd1 vssd1 vccd1 vccd1 _3424_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3544__C _4911_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3868__A1 _5773_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3355_ _3355_/A vssd1 vssd1 vccd1 vccd1 _3355_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4937__A _4937_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3286_ _3292_/A _5535_/Q vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__and2_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5025_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5085__A3 _5066_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2843__A2 _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4094__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4672__A _4672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4045__A1 _5468_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5242__B1 _4848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3288__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _5543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5789_ _5802_/CLK _5789_/D vssd1 vssd1 vccd1 vccd1 _5789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2920__A _3699_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5653__D _5653_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5008__A _5008_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4269__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4847__A _5066_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5443__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input147_A spi_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__A1 _5484_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4243__B_N _3770_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5593__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4582__A _4592_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5233__B1 _2550_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output199_A _4249_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5563__D _5563_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output366_A _3022_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2976__S _3251_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4757__A _4757_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3140_ _4335_/B _5401_/Q _3151_/S vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3380__B _3380_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5067__A3 _5066_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3071_ _5138_/C _5320_/Q _4375_/A vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__mux2_8
XFILLER_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2825__A2 _2745_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4492__A _4492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3600__S _3600_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2724__B _2724_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3973_ _4145_/A _4079_/B _3973_/C vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__and3_2
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5738__D _5738_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5712_ _5766_/CLK _5712_/D vssd1 vssd1 vccd1 vccd1 _5712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3786__B1 _3776_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2924_ _3530_/A vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5643_ _5659_/CLK _5643_/D vssd1 vssd1 vccd1 vccd1 _5643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5316__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2855_ _3711_/A _2854_/X _5486_/Q vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__3836__A _4117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2740__A _2780_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5574_ _5586_/CLK _5574_/D vssd1 vssd1 vccd1 vccd1 _5574_/Q sky130_fd_sc_hd__dfxtp_1
X_2786_ _5759_/Q _3047_/A _2658_/Y _2540_/X vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__3555__B _3565_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4525_ _4525_/A vssd1 vssd1 vccd1 vccd1 _5412_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4116__B_N _4083_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5473__D _5473_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5466__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4456_ _4891_/A _4473_/B _4456_/C vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__or3_1
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3407_ _3407_/A vssd1 vssd1 vccd1 vccd1 _3435_/S sky130_fd_sc_hd__buf_2
XFILLER_63_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4667__A _4667_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4387_ _4387_/A vssd1 vssd1 vccd1 vccd1 _5352_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3571__A _3571_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3338_ _4306_/A _5492_/Q _3441_/S vssd1 vssd1 vccd1 vccd1 _4683_/C sky130_fd_sc_hd__mux2_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__B _4425_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3290__B _5537_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _4390_/A _5528_/Q _3444_/S vssd1 vssd1 vccd1 vccd1 _4771_/C sky130_fd_sc_hd__mux2_4
XANTENNA__4266__A1 _2728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5008_/A vssd1 vssd1 vccd1 vccd1 _5635_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5648__D _5648_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3241__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3746__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2650__A _2650_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5383__D _5383_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2752__A1 _2675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3481__A _3481_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__B1 _3696_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__A2 _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4009__A1 _5781_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4009__B2 _4008_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5201__A _5201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2544__B _2544_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5558__D _5558_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5339__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5489__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2640_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__buf_4
XANTENNA__2560__A _5695_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4193__B1 _4187_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2571_ _5361_/Q _2565_/X _2570_/Y vssd1 vssd1 vccd1 vccd1 _2589_/C sky130_fd_sc_hd__o21ai_1
Xoutput306 _3531_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[31] sky130_fd_sc_hd__buf_2
Xoutput317 _3578_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput328 _3614_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[21] sky130_fd_sc_hd__buf_2
XANTENNA__2743__A1 _2698_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4310_ _4310_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__or2_1
Xoutput339 _3647_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[31] sky130_fd_sc_hd__buf_2
X_5290_ _5781_/Q _5289_/X _3993_/X _4008_/Y _5285_/X vssd1 vssd1 vccd1 vccd1 _5781_/D
+ sky130_fd_sc_hd__o221a_1
X_4241_ _3878_/A _4095_/X _5481_/Q vssd1 vssd1 vccd1 vccd1 _4241_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__4487__A _4487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3391__A _3391_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4172_ _4252_/A _4172_/B _4252_/C _4172_/D vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__and4_4
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _3123_/A _3134_/B _4487_/C vssd1 vssd1 vccd1 vccd1 _3124_/A sky130_fd_sc_hd__and3_1
XFILLER_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4248__A1 _5797_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4248__B2 _4247_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3054_ _3062_/A _3073_/B _4458_/A vssd1 vssd1 vccd1 vccd1 _3055_/A sky130_fd_sc_hd__and3_1
XFILLER_97_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4799__A2 _4780_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4934__B _4938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5111__A _5111_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5468__D _5468_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4950__A _4950_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3956_ _3956_/A1 _3954_/X _3714_/X _3955_/Y vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__a31oi_4
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4420__A1 _5369_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2907_ _2826_/X _2717_/Y _2906_/Y vssd1 vssd1 vccd1 vccd1 _2908_/D sky130_fd_sc_hd__a21oi_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _4059_/A vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__buf_4
XANTENNA__3566__A _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2982__A1 _2973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5626_ _5692_/CLK _5626_/D vssd1 vssd1 vccd1 vccd1 _5626_/Q sky130_fd_sc_hd__dfxtp_1
X_2838_ _2835_/Y _2837_/X _2864_/A vssd1 vssd1 vccd1 vccd1 _2909_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2901__C _2935_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4184__B1 _3846_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5557_ _5802_/CLK _5557_/D vssd1 vssd1 vccd1 vccd1 _5557_/Q sky130_fd_sc_hd__dfxtp_1
X_2769_ _2877_/A _2879_/A _2909_/C _2768_/Y _5556_/Q vssd1 vssd1 vccd1 vccd1 _3736_/A
+ sky130_fd_sc_hd__a41oi_4
X_4508_ _4508_/A _4526_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__and3_1
X_5488_ _5586_/CLK _5488_/D vssd1 vssd1 vccd1 vccd1 _5488_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5279__A3 _5069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4439_ _4439_/A _4439_/B _4439_/C vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__or3_1
XANTENNA__4397__A _4397_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4828__C _4988_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3732__C _3732_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5005__B _5005_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4239__B2 _3808_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2645__A _2645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3240__S _3240_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3462__A2 _2927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5021__A _5021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2670__B1 _4441_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5378__D _5378_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4860__A _5089_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5631__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3907__C _3907_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input75_A gpio_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4175__B1 _4174_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5781__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2725__A1 _2631_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3415__S _3435_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3150__A1 _5333_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output231_A _3324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output329_A _3618_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4754__B _4763_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2555__A _2809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3150__S _3162_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4473__C _4473_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4650__A1 _5472_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2661__B1 _2699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _4171_/A vssd1 vssd1 vccd1 vccd1 _4240_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__4770__A _4770_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4790_ _4801_/A _5535_/Q _4796_/C vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__and3_1
XFILLER_57_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3741_ _3720_/X _3722_/X _3733_/X _3738_/X _3740_/X vssd1 vssd1 vccd1 vccd1 _3741_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3672_ _5058_/B _2919_/A _5693_/Q vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_18_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5690_/CLK sky130_fd_sc_hd__clkbuf_16
X_5411_ _5531_/CLK _5411_/D vssd1 vssd1 vccd1 vccd1 _5411_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4166__B1 _4165_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2623_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2695_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__2716__A1 _2607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3913__B1 _3900_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5342_ _5731_/CLK _5342_/D vssd1 vssd1 vccd1 vccd1 _5342_/Q sky130_fd_sc_hd__dfxtp_1
X_2554_ _5382_/Q vssd1 vssd1 vccd1 vccd1 _2809_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5115__C1 _4883_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5273_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5751__D _5751_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3552__C _4915_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__A _4036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4224_ _4224_/A vssd1 vssd1 vccd1 vccd1 _4224_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5504__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4155_ _5790_/Q _4070_/X _4143_/X _4154_/Y vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__4945__A _4963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3106_ _3106_/A vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__clkbuf_1
X_4086_ _4081_/Y _3906_/X _4085_/Y vssd1 vssd1 vccd1 vccd1 _4086_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5654__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4680__A _4680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4988_ _4988_/A _4988_/B _4988_/C vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__and3_1
XFILLER_36_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3939_ _5462_/Q _3815_/X _3938_/X vssd1 vssd1 vccd1 vccd1 _3939_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__3296__A _3296_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2955__A1 input13/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2631__C _2929_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5609_ _5641_/CLK _5609_/D vssd1 vssd1 vccd1 vccd1 _5609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3697__C_N _3670_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3904__B1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5106__C1 _4200_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5661__D _5661_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3235__S _3235_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4558__C _4558_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3132__A1 _5330_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4855__A _5090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4880__A1 _4875_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2643__B1 _2642_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4590__A _4590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3199__A1 _5411_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3918__B _3918_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3637__C _4978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput16 cpu_adr_i[22] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 cpu_adr_i[3] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput38 cpu_dat_i[12] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 cpu_dat_i[22] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output181_A _3987_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output279_A _3454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3934__A _4141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4749__B _4763_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5527__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5571__D _5571_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3145__S _3192_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5112__A2 _4988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2984__S _3251_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4765__A _4765_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4871__A1 _4859_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5677__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_7_CLK clkbuf_leaf_7_CLK/A vssd1 vssd1 vccd1 vccd1 _5435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4911_ _4911_/A _4915_/B _4915_/C vssd1 vssd1 vccd1 vccd1 _4912_/A sky130_fd_sc_hd__and3_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4842_ _4971_/A vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__buf_4
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4773_/A _4778_/B _4778_/C vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__and3_1
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5746__D _5746_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3724_ _3998_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3547__C _4913_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4005__A _4005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2850__A_N _2846_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3655_ _3482_/A _2927_/A _4905_/C vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3844__A _4091_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2606_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__clkbuf_4
X_3586_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3601_/B sky130_fd_sc_hd__clkbuf_1
X_5325_ _5766_/CLK _5325_/D vssd1 vssd1 vccd1 vccd1 _5325_/Q sky130_fd_sc_hd__dfxtp_1
X_2537_ _2543_/A _2652_/A _5382_/Q vssd1 vssd1 vccd1 vccd1 _2573_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5481__D _5481_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2570__C1 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4170__A2_N _5684_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5256_ _5256_/A vssd1 vssd1 vccd1 vccd1 _5760_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5103__A2 _5094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4207_ _4204_/Y _4115_/X _4206_/Y vssd1 vssd1 vccd1 vccd1 _4207_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4675__A _4675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5187_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4862__A1 _4859_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4394__B _4425_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2873__B1 _5268_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4069_ _4123_/A _4069_/B vssd1 vssd1 vccd1 vccd1 _4069_/Y sky130_fd_sc_hd__nor2_8
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2626__C _2836_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2923__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5656__D _5656_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2928__A1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3050__A0 _5130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3754__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input177_A spi_rty_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4569__B _5429_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3353__A1 _5496_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4131__A_N _3999_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5391__D _5391_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A cpu_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3656__A2 _2949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4853__A1 _3925_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4853__B2 _4833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3712__C_N _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4066__C1 _4005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2536__C _2583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4751__C _4765_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5566__D _5566_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output396_A _3172_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__A1 _5644_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5030__B2 _5011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2979__S _3246_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3664__A _3664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _3440_/A vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3371_ _3407_/A vssd1 vssd1 vccd1 vccd1 _3400_/S sky130_fd_sc_hd__buf_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2552__C1 _2611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3895__A2 _4634_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5110_ _5096_/A _4837_/A _4872_/A _5268_/A _4252_/B vssd1 vssd1 vccd1 vccd1 _5690_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5650_/Q _5033_/X _5029_/X _5034_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5650_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4495__A _4495_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4844__A1 _3798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4926__C _4926_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4844__B2 _4833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3558__B _3565_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4825_ _4828_/A _5553_/Q _4988_/C vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__and3_1
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5476__D _5476_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4756_ _4756_/A _4756_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__and3_1
XANTENNA__3583__A1 _5608_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5309__C1 _5287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3707_ _4059_/A vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__buf_2
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _5493_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3574__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3638_ _3638_/A vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3569_ _4324_/A _5604_/Q _3597_/S vssd1 vssd1 vccd1 vccd1 _4930_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5308_ _5308_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5798_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5088__A1 _5081_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _2611_/B _2611_/C _4891_/X _5238_/X vssd1 vssd1 vccd1 vccd1 _5747_/D sky130_fd_sc_hd__a211o_1
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2846__B1 _5363_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2637__B _2637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4599__B1 _4584_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5260__A1 _5764_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__A0 _4392_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5386__D _5386_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5012__A1 _5636_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5372__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5012__B2 _5011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4220__C1 _4835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3484__A _3530_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4299__B _4299_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3877__A2 _5114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5079__A1 _4889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5204__A _5204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2837__B1 _2628_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output311_A _3478_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output409_A _3232_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5251__A1 _2637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3659__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5715__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2940_ _3549_/A vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__buf_2
XANTENNA__2563__A _2573_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3262__B1 _4767_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4481__C _4485_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3801__A2 _4626_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4177__A_N _4082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2871_ _5694_/Q _4968_/A _2870_/Y vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__o21ai_4
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4610_ _5448_/Q _4573_/D _3062_/A _4590_/A _4598_/X vssd1 vssd1 vccd1 vccd1 _5448_/D
+ sky130_fd_sc_hd__a221o_1
X_5590_ _5694_/CLK _5590_/D vssd1 vssd1 vccd1 vccd1 _5590_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4541_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3394__A _3394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4472_ _4472_/A vssd1 vssd1 vccd1 vccd1 _5391_/D sky130_fd_sc_hd__clkbuf_1
X_3423_ _3429_/A _3433_/B _4741_/A vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__and3_1
XANTENNA__3868__A2 _5268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3357_/A _3361_/B _4694_/C vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__and3_1
XFILLER_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3285_/A vssd1 vssd1 vccd1 vccd1 _3285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5114__A _5114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5024_ _5642_/Q _5010_/X _5806_/A _5011_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5642_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2828__B1 _2827_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4953__A _4953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5395__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5242__A1 _5266_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4045__A2 _3815_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3253__B1 _4456_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3288__B _5536_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4808_ _4821_/A _5543_/Q _4817_/C vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__and3_1
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5788_ _5798_/CLK _5788_/D vssd1 vssd1 vccd1 vccd1 _5788_/Q sky130_fd_sc_hd__dfxtp_1
X_4739_ _4749_/A _4739_/B _4739_/C vssd1 vssd1 vccd1 vccd1 _4740_/A sky130_fd_sc_hd__or3_1
XFILLER_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__S _3251_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4108__A1_N _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4284__A2 _4444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5738__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4582__B _5435_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5233__A1 _2848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3479__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3244__A0 _4297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3795__A1 _3794_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2911__A_N _2886_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2755__C1 _2611_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output261_A _3427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output359_A _3009_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3380__C _4712_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3070_ _5705_/Q input60/X _3108_/S vssd1 vssd1 vccd1 vccd1 _5138_/C sky130_fd_sc_hd__mux2_1
XFILLER_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4773__A _4773_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3235__A0 _4373_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3972_ _3817_/X _3818_/X _3972_/C _4043_/D vssd1 vssd1 vccd1 vccd1 _3973_/C sky130_fd_sc_hd__and4bb_1
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2724__C _2724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _5765_/CLK _5711_/D vssd1 vssd1 vccd1 vccd1 _5711_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3786__A1 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2923_ _3517_/A vssd1 vssd1 vccd1 vccd1 _3530_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3786__B2 _3785_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5642_ _5659_/CLK _5642_/D vssd1 vssd1 vccd1 vccd1 _5642_/Q sky130_fd_sc_hd__dfxtp_1
X_2854_ _3709_/A _3710_/A vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__or2_2
XANTENNA__5754__D _5754_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2785_ _2785_/A vssd1 vssd1 vccd1 vccd1 _3047_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2740__B _2779_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5573_ _5694_/CLK _5573_/D vssd1 vssd1 vccd1 vccd1 _5573_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3555__C _4920_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4524_ _4538_/A _4524_/B _4524_/C vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__or3_1
XANTENNA__3943__D1 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2844__B1_N _3678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4455_ _4455_/A vssd1 vssd1 vccd1 vccd1 _5385_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4948__A _5025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3852__A _4265_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3406_ _3406_/A vssd1 vssd1 vccd1 vccd1 _3406_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4386_ _4386_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__or2_1
XFILLER_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4667__B _4681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3337_ _3407_/A vssd1 vssd1 vccd1 vccd1 _3441_/S sky130_fd_sc_hd__buf_4
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3268_ _4295_/C vssd1 vssd1 vccd1 vccd1 _3268_/X sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4266__A2 _3716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5007_ _5007_/A _5130_/B _5021_/A vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__and3_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4683__A _4699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3474__B1 _5003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3199_ _4357_/B _5411_/Q _3209_/S vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__mux2_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3299__A _3303_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3746__B _3746_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2650__B _2650_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5664__D _5664_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3238__S _3246_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5410__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2752__A2 _2750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3762__A _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3701__B2 _3700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5560__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A cpu_adr_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4593__A _4593_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4662__C1 _4630_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__D1 _2806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4009__A2 _3915_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2544__C _2583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4414__C1 _4299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3002__A _3002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2841__A _2841_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__D1 _4117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__D _5574_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4193__A1 _5105_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2570_ _2761_/A _2790_/A _2567_/Y _2559_/X _2569_/X vssd1 vssd1 vccd1 vccd1 _2570_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput307 _3468_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput318 _3582_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__2987__S _3246_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2743__A2 _2640_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput329 _3618_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[22] sky130_fd_sc_hd__buf_2
XANTENNA__4768__A _4768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4240_/A _4240_/B _4240_/C _4240_/D vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__and4_2
XANTENNA__4487__B _4498_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4171_ _4171_/A vssd1 vssd1 vccd1 vccd1 _4252_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _4329_/A _5398_/Q _3146_/S vssd1 vssd1 vccd1 vccd1 _4487_/C sky130_fd_sc_hd__mux2_1
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4248__A2 _4091_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ _4304_/B _5387_/Q _3248_/S vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4934__C _4934_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4653__C1 _4645_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5749__D _5749_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5111__B _5111_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3208__A0 _5193_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _3794_/X _3919_/X _5463_/Q vssd1 vssd1 vccd1 vccd1 _3955_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_56_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4420__A2 _5238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2906_ _2829_/Y _2903_/A _2832_/Y vssd1 vssd1 vccd1 vccd1 _2906_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2751__A _5360_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5433__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3886_ _3953_/A _3886_/B _3993_/C _4026_/D vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__and4_2
XANTENNA__2982__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5625_ _5659_/CLK _5625_/D vssd1 vssd1 vccd1 vccd1 _5625_/Q sky130_fd_sc_hd__dfxtp_1
X_2837_ _2707_/A _2836_/Y _2708_/X _2628_/C _2696_/A vssd1 vssd1 vccd1 vccd1 _2837_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5484__D _5484_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4184__A1 _5685_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4184__B2 _4184_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5556_ _5589_/CLK _5556_/D vssd1 vssd1 vccd1 vccd1 _5556_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2768_ _2852_/D _2917_/B vssd1 vssd1 vccd1 vccd1 _2768_/Y sky130_fd_sc_hd__nor2_1
X_4507_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4678__A _4678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5583__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5487_ _5531_/CLK _5487_/D vssd1 vssd1 vccd1 vccd1 _5487_/Q sky130_fd_sc_hd__dfxtp_1
X_2699_ _2699_/A vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3582__A _3582_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4438_ _4438_/A vssd1 vssd1 vccd1 vccd1 _5379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3732__D _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _5346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4892__C1 _4891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5005__C _5005_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3732__A_N _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3447__A0 _4292_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2926__A _4295_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A _5302_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__D _5659_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5021__B _5641_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2670__A1 _5381_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3757__A _3757_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5394__D _5394_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3907__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4175__A1 _5476_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2725__A2 _2724_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4588__A _4588_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input68_A cpu_sel_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3492__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3438__A0 _4368_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output224_A _3309_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2836__A _2836_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4635__C1 _4632_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4754__C _4754_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5212__A _5212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5569__D _5569_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4650__A2 _4639_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2661__B2 _2672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5456__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3740_ _4005_/A vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3699_/B _3698_/A vssd1 vssd1 vccd1 vccd1 _4139_/A sky130_fd_sc_hd__nand2_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5410_ _5531_/CLK _5410_/D vssd1 vssd1 vccd1 vccd1 _5410_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4166__A1 _4059_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2622_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2736_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2716__A2 _2549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3913__A1 _5776_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2553_ _5360_/Q _2540_/X _2552_/Y vssd1 vssd1 vccd1 vccd1 _2794_/A sky130_fd_sc_hd__o21ai_1
XFILLER_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3913__B2 _3912_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5341_ _5731_/CLK _5341_/D vssd1 vssd1 vccd1 vccd1 _5341_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4498__A _4514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5115__B1 _5060_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _5769_/Q _5269_/X _3705_/X _3744_/Y _5310_/B vssd1 vssd1 vccd1 vccd1 _5769_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4223_ _4263_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4223_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__4010__B _4010_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3677__B1 _3676_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4874__C1 _4865_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4154_ _4042_/X _4146_/Y _4152_/Y _4153_/X vssd1 vssd1 vccd1 vccd1 _4154_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4945__B _4963_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3105_ _3123_/A _3105_/B _4481_/A vssd1 vssd1 vccd1 vccd1 _3106_/A sky130_fd_sc_hd__and3_1
X_4085_ _3977_/X _3978_/X _3979_/X _4084_/X _3908_/X vssd1 vssd1 vccd1 vccd1 _4085_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5122__A _5195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3036_ _3038_/A _5448_/Q vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__and2_1
XFILLER_97_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5479__D _5479_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__A _4961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4987_ _5056_/A vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3577__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ _4283_/A _4079_/B _3938_/C vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__and3_1
XFILLER_36_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3869_ _3869_/A _3869_/B vssd1 vssd1 vccd1 vccd1 _3869_/Y sky130_fd_sc_hd__nor2_8
X_5608_ _5692_/CLK _5608_/D vssd1 vssd1 vccd1 vccd1 _5608_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3701__A1_N _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__A1 _5460_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539_ _5555_/CLK _5539_/D vssd1 vssd1 vccd1 vccd1 _5539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5106__B1 _5097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5329__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3668__B1 _5485_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4880__A2 _4876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2656__A _2780_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3251__S _3251_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5032__A _5032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5479__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input122_A ksc_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__D _5389_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__B1 _4092_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__C1 _5285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2643__A1 _5378_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3918__C _3993_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput17 cpu_adr_i[23] vssd1 vssd1 vccd1 vccd1 _2734_/C sky130_fd_sc_hd__clkbuf_4
Xinput28 cpu_adr_i[4] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
Xinput39 cpu_dat_i[13] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4749__C _4749_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5207__A _5207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output341_A _3553_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3950__A _4287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4765__B _4778_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4871__A2 _4860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__A input4/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3161__S _3186_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5281__C1 _5310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4910_ _4910_/A vssd1 vssd1 vccd1 vccd1 _5596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4781__A _4781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _4836_/X _4837_/X _3774_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5558_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3397__A _3412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4772_ _4772_/A vssd1 vssd1 vccd1 vccd1 _5528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3723_ _3957_/A vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3654_ _4301_/A _5594_/Q _3654_/S vssd1 vssd1 vccd1 vccd1 _4905_/C sky130_fd_sc_hd__mux2_1
XFILLER_88_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2605_ _5362_/Q vssd1 vssd1 vccd1 vccd1 _2605_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5762__D _5762_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3585_ _3585_/A vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__clkbuf_1
X_5324_ _5765_/CLK _5324_/D vssd1 vssd1 vccd1 vccd1 _5324_/Q sky130_fd_sc_hd__dfxtp_1
X_2536_ _5768_/Q _2581_/A _2583_/A vssd1 vssd1 vccd1 vccd1 _2652_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__2570__B1 _2567_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4956__A _4956_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5255_ _5255_/A _5266_/B _5264_/C vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__and3_1
XFILLER_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5103__A3 _5087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3860__A _4082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4206_ _3763_/A _3766_/A _3768_/A _4205_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4206_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__5621__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5186_ _5200_/A _5191_/B _5186_/C vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__or3_1
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4862__A2 _4860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4137_ _4195_/A _4137_/B vssd1 vssd1 vccd1 vccd1 _4137_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3071__S _4375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2873__A1 _2776_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ _5785_/Q _3915_/X _4058_/X _4067_/Y vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__o22ai_4
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2626__D _2695_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5272__C1 _5310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5771__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3019_ _3027_/A _5440_/Q vssd1 vssd1 vccd1 vccd1 _3020_/A sky130_fd_sc_hd__and2_1
XANTENNA__4691__A _4691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3822__B1 _3821_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5024__C1 _5023_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3100__A _3100_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2928__A2 _2596_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3050__A1 _5317_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5672__D _5672_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3246__S _3246_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3889__B1 _3888_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5027__A _5043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4569__C _4665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3770__A _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4853__A2 _3926_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4066__B1 _4064_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4106__A _4123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3010__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__A2 _5010_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output291_A _3503_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output389_A _3130_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5582__D _5582_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3156__S _3192_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3370_ _3370_/A vssd1 vssd1 vccd1 vccd1 _3370_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5644__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2552__B1 _2550_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4776__A _4913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3680__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5040_ _5040_/A vssd1 vssd1 vccd1 vccd1 _5649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4844__A2 _3799_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5794__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2855__A1 _3711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__D _5757_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4824_ _5552_/Q _4803_/A _3339_/A _4804_/A _4823_/X vssd1 vssd1 vccd1 vccd1 _5552_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3558__C _4924_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4755_ _4755_/A vssd1 vssd1 vccd1 vccd1 _5520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3855__A _4846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5309__B1 _4273_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3706_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__buf_2
X_4686_ _4686_/A _4707_/B _4690_/C vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__and3_1
XANTENNA__3574__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2791__B1 _5747_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3637_ _3646_/A _3637_/B _4978_/A vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__and3_1
XANTENNA__5492__D _5492_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3066__S _3102_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3568_ _3608_/A vssd1 vssd1 vccd1 vccd1 _3597_/S sky130_fd_sc_hd__buf_2
X_5307_ _5797_/Q _5268_/D _4240_/X _4247_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5797_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4686__A _4686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3499_ _3499_/A vssd1 vssd1 vccd1 vccd1 _3499_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5088__A2 _5078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5238_ _5238_/A vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__buf_4
XFILLER_44_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _5169_/A _5178_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5170_/A sky130_fd_sc_hd__and3_1
XANTENNA__2846__A1 _2806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2637__C _2637_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5245__C1 _5238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4599__A1 _5442_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4599__B2 _4590_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5310__A _5310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5260__A2 _5234_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__A1 _5529_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5667__D _5667_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5517__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5012__A2 _5010_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4220__B1 _4218_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3765__A _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5667__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input50_A cpu_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4596__A _4611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5079__A2 _5078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2837__A1 _2707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3005__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4039__B1 _4038_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output304_A _3464_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5220__A _5220_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5251__A2 _2637_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3798__C1 _3797_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3262__A1 _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5577__D _5577_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2870_ _2861_/Y _3455_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _2870_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4540_ _4567_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__buf_6
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4471_ _4471_/A _4475_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__and3_1
X_3422_ _4357_/B _5515_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _4316_/A _5496_/Q _3441_/S vssd1 vssd1 vccd1 vccd1 _4694_/C sky130_fd_sc_hd__mux2_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3292_/A _5534_/Q vssd1 vssd1 vccd1 vccd1 _3285_/A sky130_fd_sc_hd__and2_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5023_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__buf_2
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 _2826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4953__B _4965_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5130__A _5130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5242__A2 _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3253__A1 _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5487__D _5487_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4807_ _4828_/A vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _5802_/CLK _5787_/D vssd1 vssd1 vccd1 vccd1 _5787_/Q sky130_fd_sc_hd__dfxtp_1
X_2999_ _3005_/A _5431_/Q vssd1 vssd1 vccd1 vccd1 _3000_/A sky130_fd_sc_hd__and2_1
XANTENNA__3585__A _3585_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4738_ _4738_/A vssd1 vssd1 vccd1 vccd1 _5513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2764__B1 _5748_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4669_ _4746_/A vssd1 vssd1 vccd1 vccd1 _4778_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2929__A _2929_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2648__B _2761_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4582__C _4665_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5040__A _5040_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5233__A2 _5227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3244__A1 _5384_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5397__D _5397_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3795__A2 _3716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input98_A gpio_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3495__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2755__B1 _2794_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output254_A _3406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5215__A _5223_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3180__A0 _5723_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output421_A _3253_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4773__B _4778_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4144__A_N _4075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2574__A _2574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3235__A1 _5418_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _4265_/A vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2724__D _2724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5710_ _5766_/CLK _5710_/D vssd1 vssd1 vccd1 vccd1 _5710_/Q sky130_fd_sc_hd__dfxtp_1
X_2922_ _5660_/Q vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__buf_2
XANTENNA__3786__A2 _5770_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5641_ _5641_/CLK _5641_/D vssd1 vssd1 vccd1 vccd1 _5641_/Q sky130_fd_sc_hd__dfxtp_1
X_2853_ _2853_/A _2853_/B _2853_/C vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__nand3_4
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3609__S _3636_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ _5586_/CLK _5572_/D vssd1 vssd1 vccd1 vccd1 _5572_/Q sky130_fd_sc_hd__dfxtp_1
X_2784_ _2783_/X _2671_/Y _2574_/X _2661_/Y vssd1 vssd1 vccd1 vccd1 _2787_/C sky130_fd_sc_hd__a31oi_1
XANTENNA__2740__C _2779_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2746__B1 _2745_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4523_ _4523_/A vssd1 vssd1 vccd1 vccd1 _5411_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3943__C1 _3942_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4454_ _4454_/A _4475_/B _4542_/A vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__and3_1
X_3405_ _3412_/A _3416_/B _4729_/C vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__and3_1
XANTENNA__5770__D _5770_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2749__A _2749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4425_/B sky130_fd_sc_hd__buf_4
XANTENNA__4667__C _4667_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5125__A _5125_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3336_ _3336_/A vssd1 vssd1 vccd1 vccd1 _3336_/X sky130_fd_sc_hd__clkbuf_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5362__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4964__A _4964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3329_/A vssd1 vssd1 vccd1 vccd1 _3267_/X sky130_fd_sc_hd__clkbuf_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5006_ _5006_/A vssd1 vssd1 vccd1 vccd1 _5634_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4120__C1 _4119_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3474__A1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4683__B _4688_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3198_ _5189_/A _5341_/Q _3219_/S vssd1 vssd1 vccd1 vccd1 _4357_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4162__B_N _3770_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3299__B _5541_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2985__A0 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4204__A _5582_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2737__B1 _4427_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5705__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2659__A _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5680__D _5680_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3162__A0 _5174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input152_A spi_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4662__B1 _4266_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input13_A cpu_adr_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2673__C1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4414__B1 _2600_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2544__D _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2976__A0 _5219_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2841__B _2909_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4178__C1 _4177_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4114__A _5576_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4193__A2 _3848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__C1 _3924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output371_A _3033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3953__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput308 _3472_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput319 _3585_/X vssd1 vssd1 vccd1 vccd1 ksc_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5385__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2569__A _2660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5590__D _5590_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3164__S _3209_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4487__C _4487_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4170_ _4139_/X _5684_/Q _4169_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _4172_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3121_ _5157_/C _5328_/Q _3132_/S vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__mux2_8
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3052_ _3163_/A vssd1 vssd1 vccd1 vccd1 _3248_/S sky130_fd_sc_hd__buf_2
XFILLER_83_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4653__B1 _4145_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3208__A1 _5343_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__A_N _5801_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3954_ _4128_/A vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__buf_4
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2967__B1 _4550_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2905_ _2690_/Y _5195_/A _2932_/C _2932_/D _2701_/Y vssd1 vssd1 vccd1 vccd1 _2908_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5765__D _5765_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3885_ _4057_/A vssd1 vssd1 vccd1 vccd1 _4026_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5624_ _5690_/CLK _5624_/D vssd1 vssd1 vccd1 vccd1 _5624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2836_ _2836_/A vssd1 vssd1 vccd1 vccd1 _2836_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5555_ _5555_/CLK _5555_/D vssd1 vssd1 vccd1 vccd1 _5555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4184__A2 _4986_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4959__A _4963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2767_ _2795_/A _2795_/D vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__nand2_2
XFILLER_69_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5728__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__A0 _4340_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4506_ _4971_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5486_ _5798_/CLK _5486_/D vssd1 vssd1 vccd1 vccd1 _5486_/Q sky130_fd_sc_hd__dfxtp_1
X_2698_ _2698_/A _2831_/B _2813_/C _2831_/D vssd1 vssd1 vccd1 vccd1 _2698_/Y sky130_fd_sc_hd__nand4_2
X_4437_ _4441_/A _4437_/B _4437_/C vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__and3_1
XFILLER_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4368_ _4368_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__or2_1
XANTENNA__4892__B1 _4280_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A cpu_adr_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3319_ _3325_/A _5550_/Q vssd1 vssd1 vccd1 vccd1 _3320_/A sky130_fd_sc_hd__and2_1
XANTENNA__4694__A _4699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A _4299_/B vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__and2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3447__A1 _5487_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__B _5308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__A _3163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5021__C _5039_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2670__A2 _2691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2958__A0 _5213_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5675__D _5675_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4175__A2 _4074_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3383__A0 _4333_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4100__C _4100_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3438__A1 _5520_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4635__B1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4109__A _4109_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output217_A _3296_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3013__A _3013_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2843__B1_N _5802_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2852__A _2852_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5585__D _5585_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3670_ _3670_/A1 _2867_/X _5694_/Q vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2621_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__buf_4
XANTENNA__4166__A2 _4654_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4779__A _4779_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3683__A _3683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4571__C1 _4565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5340_ _5737_/CLK _5340_/D vssd1 vssd1 vccd1 vccd1 _5340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2552_ _2848_/A _2790_/A _2550_/Y _2611_/A vssd1 vssd1 vccd1 vccd1 _2552_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__3913__A2 _3804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4498__B _4498_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4093__A1_N _3989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5115__A1 _5694_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5271_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5310_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5115__B2 _5114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3126__A0 _5714_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4222_ _5795_/Q _4091_/X _4214_/X _4221_/Y vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__o22ai_4
XANTENNA__3677__A1 _4746_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4874__B1 _4872_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4153_ _4153_/A vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4945__C _4945_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3104_ _4322_/B _5395_/Q _3151_/S vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _4082_/X _4083_/X _4084_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__and4bb_1
XFILLER_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3035_ _3035_/A vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5400__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4961__B _4965_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3858__A _4005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4986_ _4986_/A vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__buf_2
XANTENNA__3577__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3937_ _3817_/X _3818_/X _3937_/C _4043_/D vssd1 vssd1 vccd1 vccd1 _3938_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__5495__D _5495_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5550__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3868_ _5773_/Q _5268_/D _3867_/Y vssd1 vssd1 vccd1 vccd1 _3869_/B sky130_fd_sc_hd__o21ai_4
X_5607_ _5692_/CLK _5607_/D vssd1 vssd1 vccd1 vccd1 _5607_/Q sky130_fd_sc_hd__dfxtp_1
X_2819_ _2819_/A _2848_/B _2848_/C _2848_/D vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__4689__A _4689_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3799_ _4830_/B _3737_/X _5559_/Q vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__o21a_1
X_5538_ _5538_/CLK _5538_/D vssd1 vssd1 vccd1 vccd1 _5538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3904__A2 _3815_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5106__A1 _5096_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5469_ _5482_/CLK _5469_/D vssd1 vssd1 vccd1 vccd1 _5469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3668__A1 _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2937__A _2937_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2656__B _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__B1 _3993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4093__B2 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4205__A_N _4082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A ksc_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2643__A2 _2565_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A _3768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2672__A _2672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3487__B _5639_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3918__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput18 cpu_adr_i[24] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input80_A gpio_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 cpu_adr_i[5] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3356__A0 _4318_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3108__A0 _5711_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3008__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output334_A _3635_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4765__C _4765_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5223__A _5223_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5423__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2619__C1 _2574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5281__B1 _3886_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3678__A _3678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5573__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2582__A _2647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4840_ _5268_/A vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3397__B _3397_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4771_ _4771_/A _4776_/B _4771_/C vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__or3_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3722_ _4062_/A vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__buf_4
XANTENNA__4792__C1 _4783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _3482_/A _2927_/A _4903_/A vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3347__A0 _4310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2604_ _2841_/A vssd1 vssd1 vccd1 vccd1 _2909_/A sky130_fd_sc_hd__buf_2
XANTENNA__4302__A _4302_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3584_ _3594_/A _3584_/B _4938_/C vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__and3_1
X_5323_ _5766_/CLK _5323_/D vssd1 vssd1 vccd1 vccd1 _5323_/Q sky130_fd_sc_hd__dfxtp_1
X_2535_ _5767_/Q vssd1 vssd1 vccd1 vccd1 _2543_/A sky130_fd_sc_hd__inv_2
XANTENNA__2570__A1 _2761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5254_ _2711_/Y _5227_/A _2712_/Y vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__o21ai_1
X_4205_ _4082_/X _4083_/X _4205_/C _4257_/D vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__and4bb_1
XFILLER_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5185_ _5185_/A vssd1 vssd1 vccd1 vccd1 _5724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5133__A _5152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4136_ _5789_/Q _4091_/X _4127_/X _4135_/Y vssd1 vssd1 vccd1 vccd1 _4137_/B sky130_fd_sc_hd__o22ai_4
XANTENNA__2873__A2 _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4972__A _5183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4067_ _4059_/X _4647_/B _4066_/Y _4007_/X vssd1 vssd1 vccd1 vccd1 _4067_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_77_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5272__B1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3018_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3027_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3822__A1 _5456_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3588__A _3594_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5024__B1 _5806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4969_ _4990_/A _4990_/B _4969_/C vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__or3_1
XFILLER_75_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4232__D1 _4117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3338__A0 _4306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5308__A _5308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4212__A _4212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3889__A1 _3889_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5027__B _5643_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4569__D _4573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4241__B1_N _5481_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5446__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2667__A _2667_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2849__C1 _2565_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5043__A _5043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5596__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4066__A1 _3997_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5263__B1 _2668_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4066__B2 _4065_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3498__A _3504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__B _4106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3010__B _5436_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output284_A _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5218__A _5218_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3961__A _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2552__A1 _2848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4776__B _4776_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3680__B _3757_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2577__A _2785_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2855__A2 _2854_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5254__B1 _2712_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3201__A _3201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4823_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5319__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4754_ _4771_/A _4763_/B _4754_/C vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__or3_1
XFILLER_33_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3705_ _3953_/A _3705_/B _5090_/A _3792_/D vssd1 vssd1 vccd1 vccd1 _3705_/X sky130_fd_sc_hd__and4_2
XANTENNA__5309__A1 _5799_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4685_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5773__D _5773_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3347__S _3441_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5128__A _5128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2791__A1 _5261_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3574__C _4932_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3636_ _4366_/B _5623_/Q _3636_/S vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5469__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3567_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3584_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4967__A _5156_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5306_ _5306_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5796_/D sky130_fd_sc_hd__nand2_1
XANTENNA__4269__B_N _3861_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3498_ _3504_/A _5644_/Q vssd1 vssd1 vccd1 vccd1 _3499_/A sky130_fd_sc_hd__and2_1
XANTENNA__4686__B _4707_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5088__A3 _5087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5237_ _5746_/Q _5234_/X _2761_/Y _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5746_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5168_ _5168_/A vssd1 vssd1 vccd1 vccd1 _5717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2846__A2 _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4119_ _4114_/Y _4115_/X _4118_/Y vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5245__B1 _4891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4599__A2 _4589_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5310__B _5310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3111__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2950__A _3157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__A1 _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4220__B2 _4219_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5683__D _5683_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4877__A _5268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3781__A _4265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4596__B _5441_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input43_A cpu_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5079__A3 _5066_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2837__A2 _2836_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3005__B _5434_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4039__B2 _3934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3798__B1 _3725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4117__A _4117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3021__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3262__A2 _2899_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5611__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5593__D _5593_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4470_ _4470_/A vssd1 vssd1 vccd1 vccd1 _5390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3421_ _3421_/A vssd1 vssd1 vccd1 vccd1 _3421_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4787__A _4801_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5761__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3352_ _3352_/A vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__clkbuf_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__D1 _2787_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3283_ _3329_/A vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A vssd1 vssd1 vccd1 vccd1 _5641_/D sky130_fd_sc_hd__clkbuf_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2828__A2 _2717_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4953__C _4965_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5768__D _5768_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5130__B _5130_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3789__B1 _3788_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4027__A _4265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3253__A2 _2882_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3866__A _4070_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2770__A _3736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4806_ _5542_/Q _4803_/X _4798_/X _4804_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5542_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2998_ _2998_/A vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__clkbuf_1
X_5786_ _5798_/CLK _5786_/D vssd1 vssd1 vccd1 vccd1 _5786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4737_ _4737_/A _4756_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__and3_1
XANTENNA__2764__A1 _2607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4668_ _4668_/A vssd1 vssd1 vccd1 vccd1 _5486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3619_ _4355_/A _5618_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _4963_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4697__A _4697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4599_ _5442_/Q _4589_/X _4584_/X _4590_/X _4598_/X vssd1 vssd1 vccd1 vccd1 _5442_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2929__B _2929_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3106__A _3106_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2648__C _2761_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5678__D _5678_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4582__D _4596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5634__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5784__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2755__A1 _2605_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3952__B1 _3951_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3942__C _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4400__A _5238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3180__A1 input48/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5215__B _5215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output247_A _3381_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3016__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output414_A _3093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4773__C _4778_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5231__A _5231_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5588__D _5588_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3970_ _4109_/A _3970_/B _4143_/C _4240_/D vssd1 vssd1 vccd1 vccd1 _3970_/X sky130_fd_sc_hd__and4_4
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2921_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5806_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3686__A _4196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2590__A _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5640_ _5659_/CLK _5640_/D vssd1 vssd1 vccd1 vccd1 _5640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2852_ _2852_/A _2852_/B _2852_/C _2852_/D vssd1 vssd1 vccd1 vccd1 _2853_/A sky130_fd_sc_hd__nor4_2
XFILLER_73_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5571_ _5694_/CLK _5571_/D vssd1 vssd1 vccd1 vccd1 _5571_/Q sky130_fd_sc_hd__dfxtp_1
X_2783_ _2813_/C _2848_/D _2848_/B _5761_/Q vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2746__A1 _2705_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2740__D _2780_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4522_ _4522_/A _4526_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__and3_1
XANTENNA__3943__B1 _3831_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__C _4013_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4453_ _5228_/A vssd1 vssd1 vccd1 vccd1 _4475_/B sky130_fd_sc_hd__clkbuf_2
X_3404_ _4346_/A _5510_/Q _3432_/S vssd1 vssd1 vccd1 vccd1 _4729_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4310__A _4310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4384_ _4384_/A vssd1 vssd1 vccd1 vccd1 _5351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2749__B _2749_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3339_/A _4761_/A _4681_/A vssd1 vssd1 vccd1 vccd1 _3336_/A sky130_fd_sc_hd__and3_1
XANTENNA__5507__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _2895_/X _2899_/X _4769_/A vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__o21a_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _5128_/A _5005_/B _5005_/C vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__or3_1
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4120__B1 _3975_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3360__S _3441_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3197_ _5726_/Q input51/X _3228_/S vssd1 vssd1 vccd1 vccd1 _5189_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3474__A2 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4683__C _4683_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5141__A _5141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5657__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5498__D _5498_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__A _4990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3596__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2985__A1 _5426_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4187__B1 _4846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_18_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5769_ _5802_/CLK _5769_/D vssd1 vssd1 vccd1 vccd1 _5769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2737__A1 _5373_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3535__S _3564_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3162__A1 _5335_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input145_A spi_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2675__A _2675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5051__A _5051_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4662__A1 _3756_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4662__B2 _4265_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2673__B1 _2671_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4890__A _5089_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4414__A1 _5365_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2976__A1 _5354_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4198__A2_N _5686_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3937__C _3937_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2841__C _2909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4178__B1 _3768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output197_A _4223_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3925__B1 _3725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3953__B _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput309 _3474_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[5] sky130_fd_sc_hd__buf_2
XFILLER_99_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output364_A _2962_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5226__A _5226_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__A_N _4075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3120_ _5713_/Q input37/X _3168_/S vssd1 vssd1 vccd1 vccd1 _5157_/C sky130_fd_sc_hd__mux2_2
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4102__B1 _5575_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3157_/A vssd1 vssd1 vccd1 vccd1 _3163_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2585__A _2585_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3180__S _3223_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4653__A1 _5474_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2664__B1 _5756_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ _3953_/A _3953_/B _3993_/C _4026_/D vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__and4_2
XANTENNA__2967__A1 _2876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4305__A _4305_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2904_ _2677_/Y _5195_/A _2814_/Y _2779_/C vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__o211a_1
X_3884_ _3695_/X _5667_/Q _3883_/Y _3700_/X vssd1 vssd1 vccd1 vccd1 _3886_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5623_ _5659_/CLK _5623_/D vssd1 vssd1 vccd1 vccd1 _5623_/Q sky130_fd_sc_hd__dfxtp_1
X_2835_ _2806_/X _2699_/X _5358_/Q vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _5555_/CLK _5554_/D vssd1 vssd1 vccd1 vccd1 _5554_/Q sky130_fd_sc_hd__dfxtp_1
X_2766_ _5363_/Q _2696_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2795_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__4959__B _4963_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__A1 _5507_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5118__C1 _4848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4505_ _4567_/A vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5781__D _5781_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5485_ _5798_/CLK _5485_/D vssd1 vssd1 vccd1 vccd1 _5485_/Q sky130_fd_sc_hd__dfxtp_1
X_2697_ _2697_/A vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__inv_2
XANTENNA__5136__A _5136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4436_ _2817_/X _2642_/Y _4402_/X vssd1 vssd1 vccd1 vccd1 _5378_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4040__A _4199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4975__A _4975_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4367_ _4367_/A vssd1 vssd1 vccd1 vccd1 _5345_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4892__A1 _4889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3318_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3318_/X sky130_fd_sc_hd__clkbuf_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4694__B _4714_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _5314_/D sky130_fd_sc_hd__clkbuf_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _2994_/A _2882_/A _4454_/A vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3090__S _3102_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2655__B1 _2654_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5021__D _5021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2958__A1 _5351_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3080__A0 _4312_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3383__A1 _5504_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5109__C1 _4240_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5691__D _5691_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3265__S _3451_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4100__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4635__A1 _5460_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2646__B1 _5366_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4109__B _4109_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2852__B _2852_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3071__A0 _5138_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4125__A _4125_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5352__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2620_ _5359_/Q _2613_/X _2619_/Y vssd1 vssd1 vccd1 vccd1 _2864_/A sky130_fd_sc_hd__o21ai_4
XFILLER_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4571__B1 _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2551_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2611_/A sky130_fd_sc_hd__buf_4
XFILLER_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3175__S _3219_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4498__C _4498_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5270_ _5270_/A _5270_/B vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__nor2_4
XANTENNA__5115__A2 _4913_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3126__A1 input38/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4221_ _4059_/X _4658_/B _4220_/Y _3840_/X vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3677__A2 _3345_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4874__A1 _4132_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4874__B2 _4873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4152_ _4147_/X _4046_/X _3975_/X _4151_/Y vssd1 vssd1 vccd1 vccd1 _4152_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__2885__B1 _5349_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3103_ _3163_/A vssd1 vssd1 vccd1 vccd1 _3151_/S sky130_fd_sc_hd__buf_2
XFILLER_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4087__C1 _4086_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3034_ _3038_/A _5447_/Q vssd1 vssd1 vccd1 vccd1 _3035_/A sky130_fd_sc_hd__and2_1
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4961__C _4965_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5776__D _5776_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4985_ _4985_/A vssd1 vssd1 vccd1 vccd1 _5626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3577__C _4934_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3936_ _4109_/A _3936_/B _4240_/C _4240_/D vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__and4_4
XFILLER_75_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3867_ _5072_/A _3848_/X _3856_/Y _3865_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _3867_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_5606_ _5692_/CLK _5606_/D vssd1 vssd1 vccd1 vccd1 _5606_/Q sky130_fd_sc_hd__dfxtp_1
X_2818_ _5377_/Q vssd1 vssd1 vccd1 vccd1 _2818_/Y sky130_fd_sc_hd__inv_2
X_3798_ _3277_/A _3723_/X _3725_/X _3797_/X vssd1 vssd1 vccd1 vccd1 _3798_/X sky130_fd_sc_hd__o211a_1
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5537_ _5538_/CLK _5537_/D vssd1 vssd1 vccd1 vccd1 _5537_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3085__S _3132_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2749_ _2749_/A _2749_/B vssd1 vssd1 vccd1 vccd1 _2879_/A sky130_fd_sc_hd__nor2_8
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5106__A2 _4837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5468_ _5798_/CLK _5468_/D vssd1 vssd1 vccd1 vccd1 _5468_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4201__C _4201_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4419_ _2826_/X _2717_/Y _4402_/X vssd1 vssd1 vccd1 vccd1 _5368_/D sky130_fd_sc_hd__a21o_1
XFILLER_87_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5399_ _5731_/CLK _5399_/D vssd1 vssd1 vccd1 vccd1 _5399_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3668__A2 _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2937__B _2937_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2656__C _2780_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3114__A _3174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A1 _5781_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__B2 _4008_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2953__A _3047_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A ksc_ack_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5375__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5686__D _5686_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3053__A0 _4304_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3784__A _4070_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 cpu_adr_i[25] vssd1 vssd1 vccd1 vccd1 _2711_/A sky130_fd_sc_hd__buf_2
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4002__C1 _4001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3356__A1 _5497_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input73_A gpio_ack_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__C _4111_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3108__A1 input66/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3008__B _5435_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5223__B _5223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output327_A _3611_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3024__A _3024_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2619__B1 _2618_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5281__A1 _5775_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5281__B2 _3895_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5718__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2863__A _2916_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5596__D _5596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3992__A1_N _3989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3397__C _4724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4770_ _4770_/A vssd1 vssd1 vccd1 vccd1 _5527_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4792__B1 _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3721_ _3755_/A vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__buf_2
XFILLER_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3694__A _4139_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3652_ _4299_/B _5593_/Q _3652_/S vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3347__A1 _5494_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2603_ _2591_/Y _2596_/X _2916_/B vssd1 vssd1 vccd1 vccd1 _2841_/A sky130_fd_sc_hd__o21a_1
X_3583_ _4333_/A _5608_/Q _3597_/S vssd1 vssd1 vccd1 vccd1 _4938_/C sky130_fd_sc_hd__mux2_1
X_5322_ _5765_/CLK _5322_/D vssd1 vssd1 vccd1 vccd1 _5322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2570__A2 _2790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5253_ _2657_/X _2658_/Y _4565_/X _5238_/X vssd1 vssd1 vccd1 vccd1 _5759_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3633__S _3633_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4204_ _5582_/Q vssd1 vssd1 vccd1 vccd1 _4204_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5184_ _5184_/A _5202_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__and3_1
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2858__B1 _3669_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5133__B _5143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4135_ _4059_/X _4651_/B _4134_/Y _4007_/X vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4048__B_N _3833_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2873__A3 _3682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4066_ _3997_/X _4062_/X _4064_/X _4065_/X _4005_/X vssd1 vssd1 vccd1 vccd1 _4066_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__5398__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5272__A1 _5769_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3869__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3017_ _3017_/A vssd1 vssd1 vccd1 vccd1 _3017_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5272__B2 _3744_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2773__A _3331_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3822__A2 _3815_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3588__B _3601_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5024__A1 _5642_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5024__B2 _5011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _4968_/A vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__buf_2
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4232__C1 _4231_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3919_ _4110_/A vssd1 vssd1 vccd1 vccd1 _3919_/X sky130_fd_sc_hd__clkbuf_2
X_4899_ _4899_/A vssd1 vssd1 vccd1 vccd1 _5591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3338__A1 _5492_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5308__B _5308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3889__A2 _4528_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5027__C _5039_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3543__S _3564_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2849__B1 _2848_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5043__B _5651_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5248__D1 _5236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5263__A1 _2667_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4066__A2 _4062_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3779__A _4074_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2683__A _2785_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3274__B1 _4776_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3498__B _5644_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3982__D1 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output277_A _3450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3019__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2552__A2 _2790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3453__S _3453_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4776__C _4776_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A _5234_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3680__C _3682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5540__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5254__A1 _2711_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3689__A _4153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3265__A0 _4388_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2593__A _2616_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5690__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822_ _4822_/A vssd1 vssd1 vccd1 vccd1 _5551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4753_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4313__A _4313_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3704_ _4057_/A vssd1 vssd1 vccd1 vccd1 _3792_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5309__A2 _5114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _5492_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2791__A2 _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5128__B _5143_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3635_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3566_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3566_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5305_ _5795_/Q _5268_/D _4214_/X _4221_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5795_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2768__A _2852_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3497_ _3497_/A vssd1 vssd1 vccd1 vccd1 _3497_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4686__C _4690_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5144__A _5144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5236_ _5236_/A vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__buf_4
XANTENNA__3884__A1_N _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4150__D1 _4117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4983__A _4983_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5167_ _5176_/A _5167_/B _5167_/C vssd1 vssd1 vccd1 vccd1 _5168_/A sky130_fd_sc_hd__or3_1
XFILLER_44_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4118_ _3977_/X _3978_/X _3979_/X _4116_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4118_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _5096_/X _5089_/X _5090_/X _5097_/X _4109_/B vssd1 vssd1 vccd1 vccd1 _5680_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5245__A1 _5244_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3599__A _3599_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3899__A1_N _3806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3256__B1 _4763_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4049_ _3977_/X _3978_/X _3979_/X _4048_/X _3908_/X vssd1 vssd1 vccd1 vccd1 _4049_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3111__B _3134_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4220__A2 _4062_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4223__A _4263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5413__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input175_A spi_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5563__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3273__S _3453_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4596__C _4604_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5054__A _5054_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input36_A cpu_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2837__A3 _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3247__A0 _5126_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3302__A _3302_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3798__A1 _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3021__B _5441_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3862__A_N _3860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output394_A _3160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3420_ _3429_/A _3433_/B _4739_/C vssd1 vssd1 vccd1 vccd1 _3421_/A sky130_fd_sc_hd__and3_1
XFILLER_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4787__B _5533_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3351_ _3357_/A _3361_/B _4690_/A vssd1 vssd1 vccd1 vccd1 _3352_/A sky130_fd_sc_hd__and3_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__C1 _2787_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3282_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3282_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5641_/Q _5039_/C _5021_/D vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__and4_1
XFILLER_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3238__A0 _5698_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4308__A _4322_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3212__A _3212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4435__C1 _4299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5130__C _5236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3789__B2 _3700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5436__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4805_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4805_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5785_ _5802_/CLK _5785_/D vssd1 vssd1 vccd1 vccd1 _5785_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5784__D _5784_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2997_ _3005_/A _5430_/Q vssd1 vssd1 vccd1 vccd1 _2998_/A sky130_fd_sc_hd__and2_1
XFILLER_37_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5139__A _5139_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4736_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4756_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2764__A2 _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4978__A _4978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4667_ _4667_/A _4681_/B _4667_/C vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__and3_1
XANTENNA__5586__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3882__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3618_ _3618_/A vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4697__B _4707_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4598_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4598_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3549_ _3549_/A vssd1 vssd1 vccd1 vccd1 _4988_/B sky130_fd_sc_hd__buf_2
XFILLER_89_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2929__C _2929_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2648__D _2761_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3477__A0 _4396_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5219_ _5223_/A _5223_/B _5219_/C vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__or3_1
XFILLER_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3229__A0 _5202_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5694__D _5694_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2755__A2 _2540_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3952__B2 _3700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3942__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5215__C _5215_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3016__B _5439_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3468__B1 _4997_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5231__B _5266_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__A _4128_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output407_A _3227_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3032__A _3038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5459__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3967__A _3967_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2920_ _3699_/B vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__clkbuf_4
X_2851_ _2760_/Y _2903_/A _2762_/Y _2589_/B vssd1 vssd1 vccd1 vccd1 _2852_/B sky130_fd_sc_hd__o211ai_1
XFILLER_34_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5570_ _5586_/CLK _5570_/D vssd1 vssd1 vccd1 vccd1 _5570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2782_ _2782_/A _2782_/B _2782_/C _2782_/D vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__nand4_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521_ _4521_/A vssd1 vssd1 vccd1 vccd1 _5410_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3943__A1 _3829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2746__A2 _2621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4798__A _4830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4013__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4452_ _4452_/A vssd1 vssd1 vccd1 vccd1 _5384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3403_ _3403_/A vssd1 vssd1 vccd1 vccd1 _3432_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4310__B _4310_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4383_ _4396_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__and2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3334_ _4304_/B _5491_/Q _3364_/S vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__mux2_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3265_ _4388_/B _5527_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__mux2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__C1 _4630_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4120__A1 _3940_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3196_ _3196_/A vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5779__D _5779_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5141__B _5154_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4038__A _4038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4980__B _4990_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2781__A _2781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4187__A1 _4185_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5768_ _5800_/CLK _5768_/D vssd1 vssd1 vccd1 vccd1 _5768_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2737__A2 _2565_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4719_ _4724_/A _4739_/B _4719_/C vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__or3_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _5765_/CLK _5699_/D vssd1 vssd1 vccd1 vccd1 _5699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4501__A _4501_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3117__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2956__A _3144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3551__S _3564_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5601__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input138_A ksc_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5689__D _5689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4662__A2 _4667_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2673__A1 _5761_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4063__A_N _3999_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4414__A2 _4400_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3787__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5751__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2691__A _2691_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3937__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2841__D _2929_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__A1 _3763_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3925__A1 _3922_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4411__A _4573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3953__C _3993_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output357_A _3004_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3027__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4886__C1 _4883_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__A _2877_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3461__S _5033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3050_ _5130_/A _5317_/Q _3102_/S vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4102__A1 _3961_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5599__D _5599_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2585__B _2848_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2649__D1 _2569_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__A2 _4652_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2664__A1 _2593_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3697__A _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ _3695_/X _5671_/Q _3951_/Y _3700_/X vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__4810__C1 _4805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2967__A2 _2882_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2903_ _2903_/A vssd1 vssd1 vccd1 vccd1 _5195_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _3883_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5622_ _5692_/CLK _5622_/D vssd1 vssd1 vccd1 vccd1 _5622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2834_ _2902_/B _2908_/C _2834_/C _2834_/D vssd1 vssd1 vccd1 vccd1 _2842_/B sky130_fd_sc_hd__nand4_4
XFILLER_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5553_ _5555_/CLK _5553_/D vssd1 vssd1 vccd1 vccd1 _5553_/Q sky130_fd_sc_hd__dfxtp_1
X_2765_ _2585_/A _2790_/A _2764_/Y _2691_/A vssd1 vssd1 vccd1 vccd1 _2850_/B sky130_fd_sc_hd__o211ai_2
XANTENNA__3636__S _3636_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4959__C _4959_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4504_ _4504_/A vssd1 vssd1 vccd1 vccd1 _5404_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5118__B1 _5060_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4321__A _4321_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5484_ _5695_/CLK _5484_/D vssd1 vssd1 vccd1 vccd1 _5484_/Q sky130_fd_sc_hd__dfxtp_1
X_2696_ _2696_/A _2696_/B _2696_/C vssd1 vssd1 vccd1 vccd1 _2932_/D sky130_fd_sc_hd__nand3_4
XANTENNA__5136__B _5154_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4435_ _5377_/Q _5238_/A _2654_/Y _4299_/A vssd1 vssd1 vccd1 vccd1 _5377_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5624__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4366_ _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__and2_1
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4892__A2 _4890_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3317_ _3325_/A _5549_/Q vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__and2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2776__A _5268_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4297_ _4297_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__or2_1
XFILLER_80_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4694__C _4694_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5152__A _5152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _4299_/B _5385_/Q _3248_/S vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4991__A _4991_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5774__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2655__A1 _5377_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ _3179_/A vssd1 vssd1 vccd1 vccd1 _3223_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3080__A1 _5391_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3546__S _3642_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5109__B1 _5102_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2591__B1 _5364_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4868__C1 _4865_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2686__A _2686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4635__A2 _4623_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2646__A1 _2809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4109__C _4143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4406__A _4406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3310__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2852__C _2852_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3071__A1 _5320_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2661__A2_N _5376_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4020__B1 _3866_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4571__A1 _5430_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4141__A _4141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4571__B2 _4564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2550_ _2707_/A _2549_/X _5745_/Q vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__5647__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3980__A _3980_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4220_ _3824_/A _4062_/X _4218_/X _4219_/X _4835_/A vssd1 vssd1 vccd1 vccd1 _4220_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4874__A2 _4133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4151_ _4148_/Y _4115_/X _4150_/Y vssd1 vssd1 vccd1 vccd1 _4151_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5797__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2885__A1 _2700_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3191__S _3223_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3102_ _5150_/A _5325_/Q _3102_/S vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__mux2_8
X_4082_ _4082_/A vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4087__B1 _3975_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3033_ _3033_/A vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4316__A _4316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4984_ _4990_/A _4990_/B _4984_/C vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__or3_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3935_ _3932_/X _5670_/Q _3933_/Y _3934_/X vssd1 vssd1 vccd1 vccd1 _3936_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3866_ _4070_/A vssd1 vssd1 vccd1 vccd1 _3866_/X sky130_fd_sc_hd__clkbuf_4
X_5605_ _5641_/CLK _5605_/D vssd1 vssd1 vccd1 vccd1 _5605_/Q sky130_fd_sc_hd__dfxtp_1
X_2817_ _2700_/X _5266_/A _5378_/Q vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5792__D _5792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4011__B1 _3846_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3797_ _3727_/X _3729_/X _3797_/C _3978_/A vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__and4bb_1
XFILLER_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5147__A _5223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5536_ _5538_/CLK _5536_/D vssd1 vssd1 vccd1 vccd1 _5536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2748_ _2782_/B _2748_/B _2782_/D _2935_/A vssd1 vssd1 vccd1 vccd1 _2749_/B sky130_fd_sc_hd__nand4_4
XANTENNA__4986__A _4986_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5467_ _5737_/CLK _5467_/D vssd1 vssd1 vccd1 vccd1 _5467_/Q sky130_fd_sc_hd__dfxtp_1
X_2679_ _2679_/A vssd1 vssd1 vccd1 vccd1 _2813_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__3890__A _4062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5106__A3 _4872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4201__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _5367_/D sky130_fd_sc_hd__clkbuf_1
X_5398_ _5731_/CLK _5398_/D vssd1 vssd1 vccd1 vccd1 _5398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4366_/A _4349_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__and2_1
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2937__C _2937_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2656__D _2782_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A2 _5289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4226__A _4252_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3130__A _3130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3053__A1 _5387_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4002__B1 _3998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5057__A _5057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_A cpu_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4896__A _4986_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4111__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3305__A _3316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5223__C _5223_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output222_A _3260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2619__A1 _2614_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5281__A2 _5269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2863__B _2916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3040__A _3042_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3975__A _4005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3720_ _4147_/A vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__buf_4
XANTENNA__4792__A1 _5536_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4792__B2 _4782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3651_ _3482_/A _2927_/A _4901_/C vssd1 vssd1 vccd1 vccd1 _3651_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3186__S _3186_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2602_ _2759_/C vssd1 vssd1 vccd1 vccd1 _2916_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3582_ _3582_/A vssd1 vssd1 vccd1 vccd1 _3582_/X sky130_fd_sc_hd__clkbuf_1
X_5321_ _5766_/CLK _5321_/D vssd1 vssd1 vccd1 vccd1 _5321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5252_ _5758_/Q _5234_/X _2687_/Y _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5758_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4203_ _5478_/Q _4074_/X _4202_/X vssd1 vssd1 vccd1 vccd1 _4203_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2858__A1 _2845_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5183_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5133__C _5133_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4134_ _3997_/X _4062_/X _4132_/X _4133_/X _4005_/X vssd1 vssd1 vccd1 vccd1 _4134_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4213__A1_N _3806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5257__C1 _4400_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2873__A4 _3683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _3961_/X _4003_/X _5573_/Q vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5272__A2 _5269_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3016_ _3016_/A _5439_/Q vssd1 vssd1 vccd1 vccd1 _3017_/A sky130_fd_sc_hd__and2_1
XANTENNA__3869__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5787__D _5787_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3588__C _4940_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4046__A _4062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5024__A2 _5010_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4967_ _5156_/A vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4232__B1 _3768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3885__A _4057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3918_ _3953_/A _3918_/B _3993_/C _4026_/D vssd1 vssd1 vccd1 vccd1 _3918_/X sky130_fd_sc_hd__and4_2
X_4898_ _4898_/A _4915_/B _4915_/C vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__and3_1
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3849_ _3849_/A vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3096__S _3132_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3889__A3 _3714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5519_ _5641_/CLK _5519_/D vssd1 vssd1 vccd1 vccd1 _5519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5027__D _5043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2849__A1 _5745_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3125__A _3212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5043__C _5056_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5248__C1 _5235_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5342__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2964__A _3144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5263__A2 _5227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input120_A ksc_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3274__A1 _3267_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5697__D _5697_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5492__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3982__C1 _3981_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2537__B1 _5382_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3019__B _5440_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3035__A _3035_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5239__C1 _5238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2874__A _5452_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5254__A2 _5227_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3265__A1 _5527_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5400__D _5400_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4821_ _4821_/A _5551_/Q _4988_/C vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__and3_1
XFILLER_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4752_ _4752_/A vssd1 vssd1 vccd1 vccd1 _5519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3703_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__clkbuf_2
X_4683_ _4699_/A _4688_/B _4683_/C vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__or3_1
XANTENNA__5309__A3 _5069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3634_ _3646_/A _3637_/B _4976_/C vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__and3_1
XANTENNA__5128__C _5128_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3565_ _3577_/A _3565_/B _4928_/A vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__and3_1
X_5304_ _5304_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5794_/D sky130_fd_sc_hd__nand2_1
X_3496_ _3504_/A _5643_/Q vssd1 vssd1 vccd1 vccd1 _3497_/A sky130_fd_sc_hd__and2_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2768__B _2917_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5365__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5235_ _5235_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4150__C1 _4149_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5166_ _5166_/A vssd1 vssd1 vccd1 vccd1 _5716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _4117_/A vssd1 vssd1 vccd1 vccd1 _4117_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5097_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5160__A _5160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5245__A2 _2648_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _3832_/X _3833_/X _4048_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__and4bb_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3256__A1 _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3111__C _4483_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4504__A _4504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3964__C1 _3743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4223__B _4223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2959__A _3157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3554__S _3642_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5708__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3192__A0 _5186_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input168_A spi_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4596__D _4596_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput290 _3501_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input29_A cpu_adr_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5070__A _5090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3247__A1 _5315_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3798__A2 _3723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2758__B1 _2757_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output387_A _3118_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5388__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4787__C _4796_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3350_ _4312_/B _5495_/Q _3364_/S vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4380__C1 _4379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__B1 _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A _5533_/Q vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__and2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5020_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5039_/C sky130_fd_sc_hd__clkbuf_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__C1 _4131_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3238__A1 input67/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4308__B _4308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4435__B1 _2654_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3639__S _3645_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4804_ _4804_/A vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4324__A _4324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5784_ _5798_/CLK _5784_/D vssd1 vssd1 vccd1 vccd1 _5784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _3042_/A vssd1 vssd1 vccd1 vccd1 _3005_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4735_ _4971_/A vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__buf_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4666_ _4666_/A vssd1 vssd1 vccd1 vccd1 _5485_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4978__B _4997_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3882__B _5280_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3617_ _3630_/A _3620_/B _4961_/A vssd1 vssd1 vccd1 vccd1 _3618_/A sky130_fd_sc_hd__and3_1
XANTENNA__2779__A _2779_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _5441_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4697__C _4716_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5155__A _5155_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3548_ _3548_/A vssd1 vssd1 vccd1 vccd1 _3548_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2929__D _2929_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4994__A _5156_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3479_ _3517_/A vssd1 vssd1 vccd1 vccd1 _3482_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5218_ _5218_/A vssd1 vssd1 vccd1 vccd1 _5738_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3477__A1 _5635_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5149_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5709_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3403__A _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3229__A1 _5347_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2988__A0 _5225_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5530__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3792__B _3792_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5680__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2912__B1 _2911_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3468__A1 _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4409__A _4567_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3313__A _3313_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5231__C _5231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3032__B _5446_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output302_A _3525_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2979__A0 _5740_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2850_ _2846_/Y _2850_/B _2850_/C _2850_/D vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__nand4b_1
XFILLER_73_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3928__C1 _3743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2781_ _2781_/A _2781_/B vssd1 vssd1 vccd1 vccd1 _2853_/B sky130_fd_sc_hd__nor2_2
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4520_ _4538_/A _4524_/B _4520_/C vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__or3_1
XFILLER_34_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3943__A2 _3830_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4451_ _4891_/A _4473_/B _4451_/C vssd1 vssd1 vccd1 vccd1 _4452_/A sky130_fd_sc_hd__or3_1
XANTENNA__3156__A0 _5172_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3402_ _3402_/A vssd1 vssd1 vccd1 vccd1 _3402_/X sky130_fd_sc_hd__clkbuf_1
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _5350_/D sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3333_ _3453_/S vssd1 vssd1 vccd1 vccd1 _3364_/S sky130_fd_sc_hd__buf_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264_ _3453_/S vssd1 vssd1 vccd1 vccd1 _3451_/S sky130_fd_sc_hd__buf_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B1 _4186_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A _5130_/B _5021_/A vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__and3_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4319__A _4319_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4120__A2 _4046_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3195_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5403__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5141__C _5160_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4980__C _4980_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2781__B _2781_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5795__D _5795_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5553__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4054__A _4123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4187__A2 _4186_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5767_ _5767_/CLK _5767_/D vssd1 vssd1 vccd1 vccd1 _5767_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4989__A _4989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2979_ _5740_/Q input29/X _3246_/S vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__mux2_2
X_4718_ _4776_/B vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__buf_2
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5698_ _5766_/CLK _5698_/D vssd1 vssd1 vccd1 vccd1 _5698_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4651_/A _4649_/B vssd1 vssd1 vccd1 vccd1 _5471_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3117__B _3134_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2673__A2 _2577_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3787__B _5275_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input96_A gpio_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4899__A _4899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__A2 _3766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3386__A0 _4335_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3925__A2 _3723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4411__B _5102_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3953__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3138__A0 _5716_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4886__B1 _4872_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3027__B _5444_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output252_A _3398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5426__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2866__B _2879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4102__A2 _4003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2649__C1 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4139__A _4139_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3043__A _3043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__C _2848_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2664__A2 _2594_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3978__A _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5576__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2882__A _2882_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5063__B1 _5204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3697__B _3697_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _3951_/A vssd1 vssd1 vccd1 vccd1 _3951_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4810__B1 _4798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _2902_/A _2902_/B _2902_/C _2902_/D vssd1 vssd1 vccd1 vccd1 _2910_/A sky130_fd_sc_hd__nand4_1
X_3882_ _3949_/A _5280_/A vssd1 vssd1 vccd1 vccd1 _3882_/Y sky130_fd_sc_hd__nor2_8
X_5621_ _5659_/CLK _5621_/D vssd1 vssd1 vccd1 vccd1 _5621_/Q sky130_fd_sc_hd__dfxtp_1
X_2833_ _2829_/Y _2565_/X _2935_/C _2832_/Y _2935_/A vssd1 vssd1 vccd1 vccd1 _2834_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_73_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5552_ _5555_/CLK _5552_/D vssd1 vssd1 vccd1 vccd1 _5552_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4602__A _4602_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2764_ _2607_/X _2708_/A _5748_/Q vssd1 vssd1 vccd1 vccd1 _2764_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4503_ _4514_/A _4524_/B _4503_/C vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__or3_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5118__A1 _5697_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5118__B2 _5114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5483_ _5798_/CLK _5483_/D vssd1 vssd1 vccd1 vccd1 _5483_/Q sky130_fd_sc_hd__dfxtp_1
X_2695_ input14/X _2695_/B _2695_/C _2695_/D vssd1 vssd1 vccd1 vccd1 _2696_/C sky130_fd_sc_hd__nand4b_4
XANTENNA__5136__C _5236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4434_ _5376_/Q _4429_/X _4433_/X _4310_/B vssd1 vssd1 vccd1 vccd1 _5376_/D sky130_fd_sc_hd__a211o_1
XFILLER_67_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _5344_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3652__S _3652_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _3316_/A vssd1 vssd1 vccd1 vccd1 _3325_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4310_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5152__B _5167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3247_ _5126_/A _5315_/Q _4375_/A vssd1 vssd1 vccd1 vccd1 _4299_/B sky130_fd_sc_hd__mux2_8
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3837__D1 _3836_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3178_ _3178_/A vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2655__A2 _2611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4014__D1 _3331_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3368__A0 _4324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4512__A _4512_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5109__A1 _5099_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2591__A1 _2569_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5449__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4868__B1 _4856_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input150_A spi_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4030__A_N _3999_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5599__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4096__A1 _4027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2646__A2 _2750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A cpu_adr_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4109__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3310__B _5546_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2852__D _2852_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4422__A _4422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__A1 _3707_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4571__A2 _4563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3038__A _3038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2877__A _2877_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _3977_/X _3978_/X _3979_/X _4149_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4150_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_9_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2885__A2 _5266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3101_ _5710_/Q input65/X _3126_/S vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4081_ _5574_/Q vssd1 vssd1 vccd1 vccd1 _4081_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5403__D _5403_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4087__A1 _3940_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3032_ _3038_/A _5446_/Q vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__and2_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3501__A _3501_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4983_ _4983_/A vssd1 vssd1 vccd1 vccd1 _5625_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4316__B _4333_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4795__C1 _4783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3934_ _4141_/A vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__buf_2
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3865_ _3824_/X _3857_/X _4835_/A _3864_/Y vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5604_ _5692_/CLK _5604_/D vssd1 vssd1 vccd1 vccd1 _5604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2816_ _2902_/A _2902_/D _2816_/C _2816_/D vssd1 vssd1 vccd1 vccd1 _2842_/A sky130_fd_sc_hd__nand4_4
XANTENNA__4332__A _4332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4011__A1 _5674_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3796_ _3796_/A1 _4528_/A _3714_/X _3795_/Y vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__a31oi_4
XANTENNA__4011__B2 _5086_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5535_ _5538_/CLK _5535_/D vssd1 vssd1 vccd1 vccd1 _5535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2747_ _2782_/A _2779_/B _2779_/D _2782_/C vssd1 vssd1 vccd1 vccd1 _2749_/A sky130_fd_sc_hd__nand4_4
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5466_ _5798_/CLK _5466_/D vssd1 vssd1 vccd1 vccd1 _5466_/Q sky130_fd_sc_hd__dfxtp_1
X_2678_ _5266_/C _2676_/X _2677_/Y vssd1 vssd1 vccd1 vccd1 _4417_/C sky130_fd_sc_hd__o21ai_1
X_4417_ _4431_/A _4417_/B _4417_/C vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__and3_1
XANTENNA__2787__A _2787_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5397_ _5446_/CLK _5397_/D vssd1 vssd1 vccd1 vccd1 _5397_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5741__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5163__A _5163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4348_ _4378_/A vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A cpu_adr_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2937__D _2937_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4279_ _3763_/X _3766_/X _3768_/X _4278_/X _3836_/X vssd1 vssd1 vccd1 vccd1 _4279_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__5313__D _5313_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4507__A _4711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4226__B _4226_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3557__S _3564_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4002__A1 _3922_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A cpu_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2697__A _2697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2721__D1 _2672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2619__A2 _2615_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3959__C _3959_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4417__A _4431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output215_A _3291_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3321__A _3325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2863__C _2916_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3040__B _5450_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4241__A1 _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5614__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4792__A2 _4780_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3467__S _3652_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3650_ _4297_/A _5592_/Q _3654_/S vssd1 vssd1 vccd1 vccd1 _4901_/C sky130_fd_sc_hd__mux2_1
XFILLER_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2601_ _5365_/Q _2637_/A _2600_/Y vssd1 vssd1 vccd1 vccd1 _2759_/C sky130_fd_sc_hd__o21ai_4
X_3581_ _3594_/A _3584_/B _4936_/A vssd1 vssd1 vccd1 vccd1 _3582_/A sky130_fd_sc_hd__and3_1
XANTENNA__5764__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3991__A _4141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5320_ _5765_/CLK _5320_/D vssd1 vssd1 vccd1 vccd1 _5320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3752__B1 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5251_ _2637_/B _2637_/C _4891_/X _5238_/X vssd1 vssd1 vccd1 vccd1 _5757_/D sky130_fd_sc_hd__a211o_1
XFILLER_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4202_ _4254_/A _4228_/B _4202_/C vssd1 vssd1 vccd1 vccd1 _4202_/X sky130_fd_sc_hd__and3_1
X_5182_ _5182_/A vssd1 vssd1 vccd1 vccd1 _5723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2858__A2 _3664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4133_ _3735_/A _4003_/X _5577_/Q vssd1 vssd1 vccd1 vccd1 _4133_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5257__B1 _4565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4064_ _3922_/X _3958_/X _3998_/X _4063_/X vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__o211a_1
X_3015_ _3015_/A vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4327__A _4344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3231__A _3236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _5619_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4232__A1 _3763_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3917_ _3695_/X _5669_/Q _3916_/Y _3700_/X vssd1 vssd1 vccd1 vccd1 _3918_/B sky130_fd_sc_hd__o2bb2ai_1
X_4897_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4915_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5158__A _5158_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4062__A _4062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3848_ _3848_/A vssd1 vssd1 vccd1 vccd1 _3848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4997__A _4997_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3779_ _4074_/A vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__buf_4
XFILLER_101_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5518_ _5635_/CLK _5518_/D vssd1 vssd1 vccd1 vccd1 _5518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5449_ _5531_/CLK _5449_/D vssd1 vssd1 vccd1 vccd1 _5449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3406__A _3406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5802_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2849__A2 _2577_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5043__D _5043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5248__B1 _2831_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4237__A _4263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3274__A2 _3268_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3141__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5637__CLK _5641_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input113_A ksc_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5787__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5068__A _5068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3982__B1 _3979_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_CLK_A clkbuf_opt_3_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2537__A1 _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4700__A _4700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3316__A _3316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5586_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output332_A _3628_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5239__B1 _4891_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4147__A _4147_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3051__A _3157_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _5207_/A vssd1 vssd1 vccd1 vccd1 _4988_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__2890__A _3665_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4751_ _4751_/A _4756_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__and3_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3197__S _3228_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3702_ _3790_/A vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__buf_2
X_4682_ _4682_/A vssd1 vssd1 vccd1 vccd1 _5491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3633_ _4364_/A _5622_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _4976_/C sky130_fd_sc_hd__mux2_1
XFILLER_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ _4322_/B _5603_/Q _3564_/S vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5303_ _5793_/Q _5114_/X _5069_/X _4193_/Y _5287_/A vssd1 vssd1 vccd1 vccd1 _5793_/D
+ sky130_fd_sc_hd__o311a_1
X_3495_ _3517_/A vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3226__A _3236_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5234_ _5234_/A vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__buf_2
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4150__B1 _3979_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5165_ _5165_/A _5178_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__and3_1
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _4082_/X _4083_/X _4116_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _4116_/X sky130_fd_sc_hd__and4bb_1
XFILLER_99_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5798__D _5798_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5160__B _5178_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4047_ _5572_/Q vssd1 vssd1 vccd1 vccd1 _4047_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4057__A _4057_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3256__A2 _2899_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4949_ _4949_/A _4965_/B _4965_/C vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__and3_1
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3964__B1 _3963_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3959__A_N _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4520__A _4538_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3192__A1 _5340_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3136__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput280 _5805_/X vssd1 vssd1 vccd1 vccd1 gpio_stb_o sky130_fd_sc_hd__buf_2
Xoutput291 _3503_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[18] sky130_fd_sc_hd__buf_2
XFILLER_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5501__D _5501_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5765_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2758__A1 _5364_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output282_A _3458_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3972__C _3972_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4380__B1 _2885_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3046__A _3212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__A1 _4415_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3280_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__clkbuf_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5802__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4132__B1 _3998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5261__A _5261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5411__D _5411_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4435__A1 _5377_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4605__A _4605_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4803_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4324__B _4333_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5783_ _5802_/CLK _5783_/D vssd1 vssd1 vccd1 vccd1 _5783_/Q sky130_fd_sc_hd__dfxtp_1
X_2995_ _2995_/A vssd1 vssd1 vccd1 vccd1 _2995_/X sky130_fd_sc_hd__clkbuf_1
X_4734_ _4734_/A vssd1 vssd1 vccd1 vccd1 _5512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4043__C _4043_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5332__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4665_ _4837_/A _4665_/B _4665_/C _4665_/D vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__and4_1
XANTENNA__4978__C _4997_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3616_ _4353_/B _5617_/Q _3636_/S vssd1 vssd1 vccd1 vccd1 _4961_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4340__A _4344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2779__B _2779_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4596_ _4611_/A _5441_/Q _4604_/C _4596_/D vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__and4_1
XFILLER_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3547_ _3558_/A _3547_/B _4913_/C vssd1 vssd1 vccd1 vccd1 _3548_/A sky130_fd_sc_hd__and3_1
XFILLER_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5482__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3478_ _3469_/X _3470_/X _5007_/A vssd1 vssd1 vccd1 vccd1 _3478_/X sky130_fd_sc_hd__o21a_1
X_5217_ _5217_/A _5225_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__and3_1
XANTENNA__2795__A _2795_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5171__A _5223_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5148_ _5152_/A _5167_/B _5148_/C vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__or3_1
XFILLER_79_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5321__D _5321_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5079_ _4889_/X _5078_/X _5066_/X _5061_/X _3918_/B vssd1 vssd1 vccd1 vccd1 _5669_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2988__A1 _5357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4515__A _4515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3792__C _3993_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4250__A _4250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2912__A1 _2900_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A cpu_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5311__C1 _5287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3468__A2 _2927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5081__A _5081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2979__A1 input29/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4425__A _4425_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5355__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3928__B1 _3927_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2780_ _2780_/A _2780_/B _2780_/C _2780_/D vssd1 vssd1 vccd1 vccd1 _2781_/B sky130_fd_sc_hd__nand4_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3475__S _3654_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5256__A _5256_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4450_ _4558_/B vssd1 vssd1 vccd1 vccd1 _4473_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3156__A1 _5334_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3401_ _3412_/A _3416_/B _4726_/A vssd1 vssd1 vccd1 vccd1 _3402_/A sky130_fd_sc_hd__and3_1
X_4381_ _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__or2_1
XANTENNA__5406__D _5406_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3332_ _3431_/A vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__clkbuf_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__B1 _4094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3263_ _3403_/A vssd1 vssd1 vccd1 vccd1 _3453_/S sky130_fd_sc_hd__clkbuf_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4656__A1 _3756_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3504__A _3504_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B2 _4185_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__buf_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3194_ _3210_/A _3194_/B _4520_/C vssd1 vssd1 vccd1 vccd1 _3195_/A sky130_fd_sc_hd__and3_1
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4335__A _4344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4054__B _5293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766_ _5766_/CLK _5766_/D vssd1 vssd1 vccd1 vccd1 _5766_/Q sky130_fd_sc_hd__dfxtp_1
X_2978_ _2973_/X _2974_/X _4554_/C vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _5505_/D sky130_fd_sc_hd__clkbuf_1
X_5697_ _5697_/CLK _5697_/D vssd1 vssd1 vccd1 vccd1 _5697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5166__A _5166_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4070__A _4070_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4648_ _5470_/Q _4639_/X _4079_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _5470_/D sky130_fd_sc_hd__a211o_1
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5316__D _5316_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4579_ _4592_/A _5433_/Q _4665_/D _4596_/D vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__and4_1
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3117__C _4485_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3414__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5378__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3083__A0 _5707_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2830__B1 _2750_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3386__A1 _5505_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input89_A gpio_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5076__A _5097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4411__C _4411_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3138__A1 input40/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__B _5545_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4886__A1 _4244_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4886__B2 _4873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output245_A _3374_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3324__A _3324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2866__C _2866_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2649__B1 _2648_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2585__D _2848_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output412_A _3082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2855__B1_N _5486_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5063__A1 _5068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3950_ _4287_/A vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__buf_8
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4810__A1 _5544_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4810__B2 _4804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2901_ _2935_/A _2935_/B _2935_/C vssd1 vssd1 vccd1 vccd1 _2902_/C sky130_fd_sc_hd__and3_1
XANTENNA__2821__B1 _2820_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3881_ _3747_/X _5774_/Q _3877_/Y _3880_/Y vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__o22ai_4
XFILLER_91_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3994__A _3994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5620_ _5692_/CLK _5620_/D vssd1 vssd1 vccd1 vccd1 _5620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2832_ _5754_/Q _2683_/X _2831_/Y _2606_/X vssd1 vssd1 vccd1 vccd1 _2832_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_73_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5551_ _5641_/CLK _5551_/D vssd1 vssd1 vccd1 vccd1 _5551_/Q sky130_fd_sc_hd__dfxtp_1
X_2763_ _2760_/Y _2696_/A _2762_/Y vssd1 vssd1 vccd1 vccd1 _2795_/A sky130_fd_sc_hd__o21ai_2
XFILLER_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4502_ _4558_/B vssd1 vssd1 vccd1 vccd1 _4524_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5118__A2 _2927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2694_ _2607_/X _2708_/A _5755_/Q vssd1 vssd1 vccd1 vccd1 _2696_/B sky130_fd_sc_hd__o21bai_4
X_5482_ _5482_/CLK _5482_/D vssd1 vssd1 vccd1 vccd1 _5482_/Q sky130_fd_sc_hd__dfxtp_1
X_4433_ _5261_/B input20/X _2708_/X _5238_/A _2783_/X vssd1 vssd1 vccd1 vccd1 _4433_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2888__B1 _5419_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4364_ _4364_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__or2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3315_/X sky130_fd_sc_hd__clkbuf_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4295_ _4466_/A _4295_/B _4295_/C _4295_/D vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__or4_4
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _5700_/Q input69/X _3246_/S vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5152__C _5152_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3837__C1 _3835_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5520__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3177_ _3183_/A _3194_/B _4512_/A vssd1 vssd1 vccd1 vccd1 _3178_/A sky130_fd_sc_hd__and3_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3065__A0 _5704_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5670__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2812__B1 _4437_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4014__C1 _4013_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3368__A1 _5500_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4512__B _4526_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5749_ _5767_/CLK _5749_/D vssd1 vssd1 vccd1 vccd1 _5749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3409__A _3412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5109__A2 _5094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__D1 _3331_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__C _4231_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2591__A2 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4868__A1 _4064_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4868__B2 _4857_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3144__A _3144_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input143_A spi_ack_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4096__A2 _4095_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2803__B1 _2932_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4703__A _5270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output195_A _4195_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__A2 _4019_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3319__A _3325_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3038__B _5449_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output362_A _3015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5543__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3054__A _3062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3100_ _3100_/A vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _5470_/Q _4074_/X _4079_/X vssd1 vssd1 vccd1 vccd1 _4080_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__3989__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4087__A2 _4046_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3031_ _3031_/A vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2893__A _4098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5693__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4982_ _4982_/A _4997_/B _4997_/C vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__and3_1
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4244__C1 _4243_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4795__B1 _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _3933_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3864_ _3859_/Y _3828_/X _3863_/Y vssd1 vssd1 vccd1 vccd1 _3864_/Y sky130_fd_sc_hd__o21ai_1
X_5603_ _5641_/CLK _5603_/D vssd1 vssd1 vccd1 vccd1 _5603_/Q sky130_fd_sc_hd__dfxtp_1
X_2815_ _2565_/X _2677_/Y _2932_/C _2814_/Y _2932_/D vssd1 vssd1 vccd1 vccd1 _2816_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3795_ _3794_/X _3716_/X _5455_/Q vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__4011__A2 _5002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5534_ _5538_/CLK _5534_/D vssd1 vssd1 vccd1 vccd1 _5534_/Q sky130_fd_sc_hd__dfxtp_1
X_2746_ _2705_/Y _2621_/X _2745_/Y vssd1 vssd1 vccd1 vccd1 _2782_/C sky130_fd_sc_hd__o21ai_2
X_5465_ _5482_/CLK _5465_/D vssd1 vssd1 vccd1 vccd1 _5465_/Q sky130_fd_sc_hd__dfxtp_1
X_2677_ _5367_/Q vssd1 vssd1 vccd1 vccd1 _2677_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4416_ _4416_/A vssd1 vssd1 vccd1 vccd1 _5366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5396_ _5731_/CLK _5396_/D vssd1 vssd1 vccd1 vccd1 _5396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2787__B _2787_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _4347_/A vssd1 vssd1 vccd1 vccd1 _5336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4278_ _3860_/X _3861_/X _4278_/C _4278_/D vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__and4bb_1
XFILLER_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3229_ _5202_/A _5347_/Q _3229_/S vssd1 vssd1 vccd1 vccd1 _4371_/B sky130_fd_sc_hd__mux2_8
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__C1 _4153_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4226__C _4252_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4523__A _4523_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5416__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4002__A2 _3958_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5566__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3573__S _3600_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5504__D _5504_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2721__C1 _2699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3602__A _3602_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3959__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4417__B _4417_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2863__D _2929_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3321__B _5551_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output208_A _3914_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4241__A2 _4095_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3049__A _3174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2600_ _2622_/A _2600_/B _2600_/C vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__nand3_1
X_3580_ _4331_/B _5607_/Q _3600_/S vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3752__A1 _4147_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3752__B2 _3662_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5264__A _5264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5250_ _2665_/B _2665_/C _5242_/Y vssd1 vssd1 vccd1 vccd1 _5756_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4201_ _4075_/X _4076_/X _4201_/C _4201_/D vssd1 vssd1 vccd1 vccd1 _4202_/C sky130_fd_sc_hd__and4bb_1
XFILLER_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3789__A1_N _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5181_ _5200_/A _5191_/B _5181_/C vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__or3_1
XANTENNA__5414__D _5414_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4132_ _4098_/X _3958_/A _3998_/X _4131_/X vssd1 vssd1 vccd1 vccd1 _4132_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5257__A1 _2783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__A _4611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4063_ _3999_/X _4000_/X _4063_/C _4063_/D vssd1 vssd1 vccd1 vccd1 _4063_/X sky130_fd_sc_hd__and4bb_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3512__A _3512_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3014_ _3016_/A _5438_/Q vssd1 vssd1 vccd1 vccd1 _3015_/A sky130_fd_sc_hd__and2_1
XFILLER_42_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4327__B _4327_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3231__B _4542_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5439__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _4965_/A _4965_/B _4965_/C vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__and3_1
XANTENNA__4232__A2 _3766_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _3916_/A vssd1 vssd1 vccd1 vccd1 _3916_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4343__A _4343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4896_ _4986_/A vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5589__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3847_ _5665_/Q _4986_/A _3846_/X _3847_/B2 vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__a22oi_4
XFILLER_14_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4997__B _4997_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3778_ _2561_/Y _3157_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__a21o_1
X_5517_ _5641_/CLK _5517_/D vssd1 vssd1 vccd1 vccd1 _5517_/Q sky130_fd_sc_hd__dfxtp_1
X_2729_ _4617_/A vssd1 vssd1 vccd1 vccd1 _5807_/A sky130_fd_sc_hd__buf_2
XANTENNA__2798__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5174__A _5174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5448_ _5531_/CLK _5448_/D vssd1 vssd1 vccd1 vccd1 _5448_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5324__D _5324_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5379_ _5695_/CLK _5379_/D vssd1 vssd1 vccd1 vccd1 _5379_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2703__C1 _2702_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5248__A1 _5754_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3259__A0 _4383_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4518__A _4518_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4237__B _5306_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3141__B _3165_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4208__C1 _4207_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A gpio_err_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3982__A1 _3977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input71_A cpu_stb_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2537__A2 _2652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5084__A _5102_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5239__A1 _2611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output325_A _3607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4428__A _4428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3332__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4043__A_N _3817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3422__A0 _4357_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4750_ _4750_/A vssd1 vssd1 vccd1 vccd1 _5518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _3695_/X _5661_/Q _3696_/Y _3700_/X vssd1 vssd1 vccd1 vccd1 _3705_/B sky130_fd_sc_hd__o2bb2ai_1
X_4681_ _4681_/A _4681_/B _4690_/C vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__and3_1
XANTENNA__5409__D _5409_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3632_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3563_ _3563_/A vssd1 vssd1 vccd1 vccd1 _3563_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3507__A _3515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2933__C1 _2932_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5302_ _5302_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5792_/D sky130_fd_sc_hd__nand2_1
X_3494_ _3494_/A vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3226__B _4542_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5233_ _2848_/A _5227_/X _2550_/Y _5228_/X _4377_/X vssd1 vssd1 vccd1 vccd1 _5745_/D
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4150__A1 _3977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5164_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5184_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4115_ _4115_/A vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4338__A _4338_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5095_ _5081_/X _5094_/X _5087_/X _5084_/X _4094_/B vssd1 vssd1 vccd1 vccd1 _5679_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5160__C _5160_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4046_ _4062_/A vssd1 vssd1 vccd1 vccd1 _4046_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3661__B1 _2800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5169__A _5169_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4073__A _4109_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4948_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4965_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4610__C1 _4598_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3964__A1 _3887_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5319__D _5319_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4879_ _4163_/X _4164_/X _4872_/X _4873_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _5579_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4801__A _4801_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4520__B _4524_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3417__A _3417_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput270 _3352_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput281 _2915_/X vssd1 vssd1 vccd1 vccd1 gpio_we_o sky130_fd_sc_hd__buf_2
Xoutput292 _3505_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[19] sky130_fd_sc_hd__buf_2
XANTENNA__5604__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3152__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2991__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5754__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3652__A0 _4299_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3404__A0 _4346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2658__A_N input18/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2758__A2 _2611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3955__A1 _3794_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5807__A _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4711__A _4711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output275_A _3370_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3972__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3327__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4380__A1 _4377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__A2 _4415_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A1 _4098_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5261__B _5261_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2694__A1 _2607_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3062__A _3062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4084__B_N _4083_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4435__A2 _5238_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5093__C1 _4073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3997__A _4147_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _5541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5782_ _5800_/CLK _5782_/D vssd1 vssd1 vccd1 vccd1 _5782_/Q sky130_fd_sc_hd__dfxtp_1
X_2994_ _2994_/A _5429_/Q vssd1 vssd1 vccd1 vccd1 _2995_/A sky130_fd_sc_hd__and2_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4733_ _4749_/A _4739_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__or3_1
XFILLER_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4043__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4621__A _4621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4664_ _4664_/A vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__buf_6
XFILLER_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3615_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__4340__B _4340_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3237__A _3237_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2779__C _2779_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3546_ _4310_/A _5598_/Q _3642_/S vssd1 vssd1 vccd1 vccd1 _4913_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5627__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3477_ _4396_/B _5635_/Q _3652_/S vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4659__C1 _4621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5216_ _5216_/A vssd1 vssd1 vccd1 vccd1 _5737_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2795__B _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5777__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5147_ _5223_/B vssd1 vssd1 vccd1 vccd1 _5167_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5602__D _5602_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5094_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_15_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4029_ _4029_/A1 _3954_/X _3994_/X _4028_/Y vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__a31oi_4
XFILLER_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3700__A _4141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4531__A _4711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__D _3792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3147__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input173_A spi_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2912__A2 _2910_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5311__B1 _3685_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A cpu_cyc_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5512__D _5512_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4706__A _4706_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3610__A _3613_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__D1 _2935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4425__B _4425_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4144__C _4144_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__A1 _3887_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output392_A _3148_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4050__B1 _4049_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4441__A _4441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3400_ _4344_/B _5509_/Q _3400_/S vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4231__A_N _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4380_ _4377_/X _5208_/A _2885_/X _4379_/X vssd1 vssd1 vccd1 vccd1 _5349_/D sky130_fd_sc_hd__o211a_1
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3331_ _3331_/A vssd1 vssd1 vccd1 vccd1 _3431_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2896__A _2909_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__A1 _5787_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__B2 _4104_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3262_ _2895_/X _2899_/X _4767_/C vssd1 vssd1 vccd1 vccd1 _3262_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3504__B _5647_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5130_/B sky130_fd_sc_hd__buf_8
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4656__A2 _4667_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193_ _4355_/A _5410_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _4520_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5422__D _5422_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3864__B1 _3863_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3616__A0 _4353_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4616__A _5207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3520__A _3526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4813__C1 _4805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4335__B _4335_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ _5765_/CLK _5765_/D vssd1 vssd1 vccd1 vccd1 _5765_/Q sky130_fd_sc_hd__dfxtp_1
X_2977_ _4390_/A _5424_/Q _3252_/S vssd1 vssd1 vccd1 vccd1 _4554_/C sky130_fd_sc_hd__mux2_1
X_4716_ _4716_/A _4731_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__and3_1
XANTENNA__4351__A _4351_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5696_ _5798_/CLK _5696_/D vssd1 vssd1 vccd1 vccd1 _5696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4647_ _4651_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _5469_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4578_ _4600_/A vssd1 vssd1 vccd1 vccd1 _4596_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3529_ _3529_/A vssd1 vssd1 vccd1 vccd1 _3529_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5182__A _5182_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5332__D _5332_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4526__A _4526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3430__A _3430_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3083__A1 input62/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2815__D1 _2932_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4280__B1 _4279_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2830__A1 _5374_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2830__B2 _2675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4032__B1 _5571_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3576__S _3597_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5507__D _5507_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4886__A2 _4245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5296__C1 _5285_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2866__D _2866_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2649__A1 _5751_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output238_A _3272_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5322__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output405_A _3217_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3340__A _3340_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5063__A2 _4664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4271__B1 _4270_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4810__A2 _4803_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2900_ _5523_/Q vssd1 vssd1 vccd1 vccd1 _2900_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2821__A1 _2818_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3880_ _3707_/X _3879_/Y _5289_/A vssd1 vssd1 vccd1 vccd1 _3880_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5472__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4072__A2_N _5678_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2831_ _2831_/A _2831_/B _2848_/C _2831_/D vssd1 vssd1 vccd1 vccd1 _2831_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__5267__A _5267_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5550_ _5555_/CLK _5550_/D vssd1 vssd1 vccd1 vccd1 _5550_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4171__A _4171_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2762_ _5746_/Q _2785_/A _2761_/Y _2704_/A _2806_/A vssd1 vssd1 vccd1 vccd1 _2762_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4501_ _4501_/A vssd1 vssd1 vccd1 vccd1 _5403_/D sky130_fd_sc_hd__clkbuf_1
X_5481_ _5482_/CLK _5481_/D vssd1 vssd1 vccd1 vccd1 _5481_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5417__D _5417_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2693_ _2675_/A _2750_/A _2692_/Y vssd1 vssd1 vccd1 vccd1 _2932_/C sky130_fd_sc_hd__o21bai_4
X_4432_ _4432_/A vssd1 vssd1 vccd1 vccd1 _5375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _5343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2888__A1 _2631_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3515__A _3515_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _3314_/A _5548_/Q vssd1 vssd1 vccd1 vccd1 _3315_/A sky130_fd_sc_hd__and2_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ input1/X vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__clkinv_2
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _2994_/A _2882_/A _4451_/C vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__o21a_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__B1 _3831_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3176_ _4349_/B _5407_/Q _3209_/S vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4346__A _4346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3065__A1 input57/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4262__B1 _4252_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2812__A1 _4427_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2812__B2 _4437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3396__S _3396_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__B1 _3768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5177__A _5177_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4081__A _5574_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5748_ _5767_/CLK _5748_/D vssd1 vssd1 vccd1 vccd1 _5748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4512__C _4512_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3409__B _3416_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5327__D _5327_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5679_ _5697_/CLK _5679_/D vssd1 vssd1 vccd1 vccd1 _5679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5109__A3 _5066_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__D _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4868__A2 _4065_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5345__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input136_A ksc_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4256__A _5586_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3160__A _3160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5495__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2803__A1 _2632_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5087__A _5087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2567__B1 _5746_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3319__B _5550_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output188_A _4106_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output355_A _3000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3335__A _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3054__B _3073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3030_ _3038_/A _5445_/Q vssd1 vssd1 vccd1 vccd1 _3031_/A sky130_fd_sc_hd__and2_1
Xinput170 spi_dat_i[4] vssd1 vssd1 vccd1 vccd1 _3851_/D sky130_fd_sc_hd__buf_2
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5700__D _5700_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _5624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4244__B1 _4781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4795__A1 _5538_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3932_ _4139_/A vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__buf_2
XANTENNA__4795__B2 _4782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _3763_/X _3766_/X _3768_/X _3862_/X _3836_/X vssd1 vssd1 vccd1 vccd1 _3863_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5602_ _5692_/CLK _5602_/D vssd1 vssd1 vccd1 vccd1 _5602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2814_ _5752_/Q _2683_/X _2813_/Y _2606_/X vssd1 vssd1 vccd1 vccd1 _2814_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3794_ _4265_/A vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2558__B1 _2544_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5533_ _5538_/CLK _5533_/D vssd1 vssd1 vccd1 vccd1 _5533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2745_ _5261_/C _2615_/X _2709_/Y _2574_/A vssd1 vssd1 vccd1 vccd1 _2745_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5464_ _5798_/CLK _5464_/D vssd1 vssd1 vccd1 vccd1 _5464_/Q sky130_fd_sc_hd__dfxtp_1
X_2676_ _2750_/A vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5368__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4415_ _4415_/A _4415_/B _4439_/C vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__or3_1
X_5395_ _5731_/CLK _5395_/D vssd1 vssd1 vccd1 vccd1 _5395_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2787__C _2787_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4180__C1 _4179_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4346_ _4346_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__or2_1
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2730__B1 _5366_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4277_ _5588_/Q vssd1 vssd1 vccd1 vccd1 _4277_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3228_ _5732_/Q input58/X _3228_/S vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4076__A _4076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3159_ _3183_/A _3165_/B _4503_/C vssd1 vssd1 vccd1 vccd1 _3160_/A sky130_fd_sc_hd__and3_1
XANTENNA__5610__D _5610_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4235__B1 _4234_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4226__D _4664_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4804__A _4804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2721__B1 _2720_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2994__A _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5520__D _5520_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_3_1_CLK_A clkbuf_opt_3_1_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4417__C _4417_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4714__A _4724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__C1 _3946_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5510__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3752__A2 _4062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5264__B _5266_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4200_ _4252_/A _4200_/B _4252_/C _4664_/A vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__and4_4
XFILLER_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5660__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2712__B1 _5760_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4131_ _3999_/X _4000_/X _4131_/C _4243_/D vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__and4bb_1
XFILLER_42_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5280__A _5280_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5257__A2 _2671_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4062_ _4062_/A vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__buf_4
XFILLER_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__B _5447_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3013_ _3013_/A vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5430__D _5430_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3231__C _4536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4964_ _4964_/A vssd1 vssd1 vccd1 vccd1 _5618_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4624__A _4645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3915_ _4091_/A vssd1 vssd1 vccd1 vccd1 _3915_/X sky130_fd_sc_hd__buf_4
X_4895_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3846_ _3846_/A vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__buf_4
XFILLER_53_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3777_ _4057_/A vssd1 vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__buf_6
XFILLER_101_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4997__C _4997_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2728_ _2728_/A vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__clkbuf_4
X_5516_ _5589_/CLK _5516_/D vssd1 vssd1 vccd1 vccd1 _5516_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2798__B _3660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2951__A0 _4381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5174__B _5178_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5447_ _5531_/CLK _5447_/D vssd1 vssd1 vccd1 vccd1 _5447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5605__D _5605_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2659_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2699_/A sky130_fd_sc_hd__buf_4
XFILLER_82_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5378_ _5695_/CLK _5378_/D vssd1 vssd1 vccd1 vccd1 _5378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2703__B1 _2689_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4329_ _4329_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__or2_1
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5190__A _5190_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5248__A2 _5234_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3703__A _4199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3259__A1 _5525_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5340__D _5340_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3141__C _4496_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4208__B1 _3758_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4534__A _4538_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5533__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3982__A2 _3978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5683__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2942__B1 _3547_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input64_A cpu_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5515__D _5515_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__A _4724_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3613__A _3613_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5239__A2 _2611_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output220_A _3302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output318_A _3582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3670__A1 _3670_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4444__A _4444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3422__A1 _5515_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _4141_/A vssd1 vssd1 vccd1 vccd1 _3700_/X sky130_fd_sc_hd__clkbuf_2
X_4680_ _4680_/A vssd1 vssd1 vccd1 vccd1 _5490_/D sky130_fd_sc_hd__clkbuf_1
X_3631_ _3631_/A vssd1 vssd1 vccd1 vccd1 _3631_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2899__A _2899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5275__A _5275_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3186__A0 _5724_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3562_ _3577_/A _3565_/B _4926_/C vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__and3_1
XANTENNA__2933__B1 _2689_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5301_ _5791_/Q _5268_/D _4159_/X _4166_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5791_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3507__B _5648_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3493_ _3493_/A _5642_/Q vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__and2_1
XANTENNA__5425__D _5425_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5232_ _5232_/A vssd1 vssd1 vccd1 vccd1 _5744_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4135__C1 _4007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3226__C _4534_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4150__A2 _3978_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5163_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3523__A _3523_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5406__CLK _5731_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4114_ _5576_/Q vssd1 vssd1 vccd1 vccd1 _4114_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _5094_/A vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4338__B _4355_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4045_ _5468_/Q _3815_/X _4044_/X vssd1 vssd1 vccd1 vccd1 _4045_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3110__A0 _4324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3661__A1 _3980_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5556__CLK _5589_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4354__A _4354_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5169__B _5178_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4947_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4073__B _4073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4610__B1 _3062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3964__A2 _4638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4878_ _4875_/X _4876_/X _4151_/Y _4877_/X vssd1 vssd1 vccd1 vccd1 _5578_/D sky130_fd_sc_hd__a211o_1
XANTENNA__4801__B _5541_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3829_ _3977_/A vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5185__A _5185_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2602__A _2759_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4520__C _4520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5335__D _5335_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput260 _3424_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput271 _3355_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput282 _3458_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput293 _3462_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__4529__A _4538_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2688__C1 _2574_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3433__A _3445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3152__B _3165_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3101__A0 _5710_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3652__A1 _5593_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3404__A1 _5510_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3955__A2 _3919_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3168__A0 _5721_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3608__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2915__B1 _4761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3327__B _5554_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4380__A2 _5208_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3873__B_N _3770_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output268_A _3446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5429__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A2 _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4439__A _4439_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3343__A _3357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5261__C _5261_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2694__A2 _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3062__B _3073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5579__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5093__B1 _5076_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4174__A _4254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2851__C1 _2589_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4801_ _4801_/A _5541_/Q _4817_/C vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__and3_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ _2993_/A vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__clkbuf_1
X_5781_ _5802_/CLK _5781_/D vssd1 vssd1 vccd1 vccd1 _5781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4732_ _4732_/A vssd1 vssd1 vccd1 vccd1 _5511_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4902__A _4902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4663_ _5484_/Q _4542_/A _4283_/X _4621_/A vssd1 vssd1 vccd1 vccd1 _5484_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3518__A _3526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3614_ _3614_/A vssd1 vssd1 vccd1 vccd1 _3614_/X sky130_fd_sc_hd__clkbuf_1
X_4594_ _5440_/Q _4589_/X _4584_/X _4590_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _5440_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2906__B1 _2832_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2779__D _2779_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3545_ _3545_/A vssd1 vssd1 vccd1 vccd1 _3545_/X sky130_fd_sc_hd__clkbuf_1
X_3476_ _3469_/X _3470_/X _5005_/C vssd1 vssd1 vccd1 vccd1 _3476_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4659__B1 _4228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5215_ _5223_/A _5215_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__or3_1
XANTENNA__4349__A _4366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2795__C _2864_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3867__D1 _3866_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5146_ _5146_/A vssd1 vssd1 vccd1 vccd1 _5708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5077_ _5075_/X _4890_/X _5070_/X _5076_/X _3900_/B vssd1 vssd1 vccd1 vccd1 _5668_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4028_ _4027_/X _3919_/X _5467_/Q vssd1 vssd1 vccd1 vccd1 _4028_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4812__A _4812_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3147__B _3165_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input166_A spi_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5311__A1 _5801_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5721__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3163__A _3163_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input27_A cpu_adr_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3610__B _3620_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__C1 _2832_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3102__S _3102_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3389__A0 _4338_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4144__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4722__A _4722_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__A2 _4636_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4050__A1 _4047_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output385_A _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4441__B _4441_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3561__A0 _4320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3330_ _3330_/A vssd1 vssd1 vccd1 vccd1 _3330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2896__B _2909_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _4386_/A _5526_/Q _3444_/S vssd1 vssd1 vccd1 vccd1 _4767_/C sky130_fd_sc_hd__mux2_4
XANTENNA__4105__A2 _4091_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5703__D _5703_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4169__A _4169_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3073__A _3092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A vssd1 vssd1 vccd1 vccd1 _5632_/D sky130_fd_sc_hd__clkbuf_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3192_ _5186_/C _5340_/Q _3192_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_8
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3864__A1 _3859_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3616__A1 _5617_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4813__B1 _4798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3520__B _5654_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4577__C1 _4576_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4632__A _4645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5764_ _5767_/CLK _5764_/D vssd1 vssd1 vccd1 vccd1 _5764_/Q sky130_fd_sc_hd__dfxtp_2
X_2976_ _5219_/C _5354_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__mux2_8
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _5504_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4351__B _4355_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5695_ _5695_/CLK _5695_/D vssd1 vssd1 vccd1 vccd1 _5695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4646_ _5468_/Q _4639_/X _4044_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _5468_/D sky130_fd_sc_hd__a211o_1
XFILLER_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4577_ _5432_/Q _4563_/X _5807_/A _4564_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _5432_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5744__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3528_ _3530_/A _5658_/Q vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__and2_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3459_ _4289_/D vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4079__A _4145_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5613__D _5613_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2648__A_N input9/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5129_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5701_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4807__A _4828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3711__A _3711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4526__B _4526_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2815__C1 _2814_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4280__A1 _4277_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2830__A2 _5376_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4542__A _4542_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4032__A1 _3961_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2997__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3543__A0 _4308_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5523__D _5523_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5296__B1 _4094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2649__A2 _2577_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4717__A _4717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3621__A _3621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output300_A _3521_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5063__A3 _4252_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4271__A1 _4268_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5617__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2821__A2 _2540_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2830_ _5374_/Q _5376_/Q _2750_/A _2675_/A vssd1 vssd1 vccd1 vccd1 _2935_/C sky130_fd_sc_hd__o22ai_2
XANTENNA__4452__A _4452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2761_ _2761_/A _2761_/B _2761_/C _2761_/D vssd1 vssd1 vccd1 vccd1 _2761_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3068__A _3092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5767__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4500_ _4500_/A _4500_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__and3_1
X_5480_ _5482_/CLK _5480_/D vssd1 vssd1 vccd1 vccd1 _5480_/Q sky130_fd_sc_hd__dfxtp_1
X_2692_ _5370_/Q vssd1 vssd1 vccd1 vccd1 _2692_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_14_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4431_ _4431_/A _4431_/B _4431_/C vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__and3_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2700__A _2806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4362_ _4366_/A _4362_/B vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__and2_1
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2888__A2 _2724_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3515__B _5652_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3313_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3313_/X sky130_fd_sc_hd__clkbuf_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5433__D _5433_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4293_/A vssd1 vssd1 vccd1 vccd1 _5313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3244_ _4297_/A _5384_/Q _3252_/S vssd1 vssd1 vccd1 vccd1 _4451_/C sky130_fd_sc_hd__mux2_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__A1 _3829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _5178_/A _5337_/Q _3219_/S vssd1 vssd1 vccd1 vccd1 _4349_/B sky130_fd_sc_hd__mux2_8
XFILLER_41_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3531__A _3531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4346__B _4355_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4262__A1 _5798_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4262__B2 _4261_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2812__A2 _4427_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4362__A _4366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__A1 _3763_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5747_ _5767_/CLK _5747_/D vssd1 vssd1 vccd1 vccd1 _5747_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5608__D _5608_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2959_ _3157_/A vssd1 vssd1 vccd1 vccd1 _3252_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3773__B1 _3768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3409__C _4731_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5678_ _5690_/CLK _5678_/D vssd1 vssd1 vccd1 vccd1 _5678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4629_ _5228_/A vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5193__A _5193_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3706__A _4199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2610__A _2610_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2733__D1 _2787_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5343__D _5343_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4537__A _4537_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input129_A ksc_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4789__C1 _4783_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3587__S _3600_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2803__A2 _2565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input94_A gpio_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5518__D _5518_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2567__A1 _2707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3335__B _4761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output250_A _3391_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output348_A _3651_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3054__C _4458_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4447__A _4466_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput160 spi_dat_i[24] vssd1 vssd1 vccd1 vccd1 _4185_/D sky130_fd_sc_hd__clkbuf_1
Xinput171 spi_dat_i[5] vssd1 vssd1 vccd1 vccd1 _3878_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__3351__A _3357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4980_ _4990_/A _4990_/B _4980_/C vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__or3_1
XANTENNA__4244__A1 _4098_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _4138_/A vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4795__A2 _4780_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5278__A _5299_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3862_ _3860_/X _3861_/X _3862_/C _4278_/D vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__and4bb_1
X_5601_ _5641_/CLK _5601_/D vssd1 vssd1 vccd1 vccd1 _5601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2813_ _2813_/A _2831_/B _2813_/C _2831_/D vssd1 vssd1 vccd1 vccd1 _2813_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__5428__D _5428_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3793_ _3849_/A vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2558__A1 _5261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5532_ _5538_/CLK _5532_/D vssd1 vssd1 vccd1 vccd1 _5532_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4910__A _4910_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2744_ _5379_/Q _2613_/X _4437_/B vssd1 vssd1 vccd1 vccd1 _2779_/D sky130_fd_sc_hd__o21ai_4
XFILLER_34_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2675_ _2675_/A vssd1 vssd1 vccd1 vccd1 _5266_/C sky130_fd_sc_hd__buf_2
X_5463_ _5741_/CLK _5463_/D vssd1 vssd1 vccd1 vccd1 _5463_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3526__A _3526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _5365_/Q _4400_/X _2600_/Y _4299_/A vssd1 vssd1 vccd1 vccd1 _5365_/D sky130_fd_sc_hd__o211a_1
X_5394_ _5731_/CLK _5394_/D vssd1 vssd1 vccd1 vccd1 _5394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2787__D _2935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4180__B1 _3758_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _5335_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4225__A1_N _4139_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2730__A1 _2809_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _5692_/Q _5002_/A _3846_/X _5112_/B2 vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_41_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3227_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3227_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4357__A _4366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3158_ _4342_/A _5404_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _4503_/C sky130_fd_sc_hd__mux2_1
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _5708_/Q input63/X _3126_/S vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4235__A1 _3792_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5188__A _5212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2605__A _5362_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__A _4092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5338__D _5338_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4820__A _5207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A _3445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_23_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5767_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2721__A1 _2831_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5462__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2994__B _5429_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5801__D _5801_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3171__A _3183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4714__B _4714_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__B1 _3984_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3110__S _3146_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output298_A _3516_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4730__A _4730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4024__A2_N _5675_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3346__A _3445_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5264__C _5264_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_14_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5555_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2712__A1 _2607_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4130_ _4130_/A1 _4449_/A _3994_/X _4129_/Y vssd1 vssd1 vccd1 vccd1 _4651_/B sky130_fd_sc_hd__a31oi_4
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4039__A2_N _5676_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5280__B _5284_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4061_ _4061_/A1 _3954_/X _3994_/X _4060_/Y vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__a31oi_4
XFILLER_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__A _3092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5711__D _5711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4608__C _5017_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3012_ _3016_/A _5437_/Q vssd1 vssd1 vccd1 vccd1 _3013_/A sky130_fd_sc_hd__and2_1
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4905__A _4913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4963_ _4963_/A _4963_/B _4963_/C vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__or3_1
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3914_ _3949_/A _5282_/A vssd1 vssd1 vccd1 vccd1 _3914_/Y sky130_fd_sc_hd__nor2_8
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4894_ _5590_/Q _4688_/B _4872_/X _4873_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _5590_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5335__CLK _5741_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3845_ _3989_/A vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3776_ _3751_/Y _5114_/A _3775_/Y vssd1 vssd1 vccd1 vccd1 _3776_/Y sky130_fd_sc_hd__o21ai_2
X_5515_ _5635_/CLK _5515_/D vssd1 vssd1 vccd1 vccd1 _5515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2727_ _3849_/A vssd1 vssd1 vccd1 vccd1 _2728_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2951__A1 _5420_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5174__C _5184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput420 _3249_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[2] sky130_fd_sc_hd__buf_2
X_5446_ _5446_/CLK _5446_/D vssd1 vssd1 vccd1 vccd1 _5446_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5485__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2658_ input18/X _2695_/B _2695_/C _2695_/D vssd1 vssd1 vccd1 vccd1 _2658_/Y sky130_fd_sc_hd__nand4b_4
X_5377_ _5695_/CLK _5377_/D vssd1 vssd1 vccd1 vccd1 _5377_/Q sky130_fd_sc_hd__dfxtp_1
X_2589_ _2794_/A _2589_/B _2589_/C _4411_/C vssd1 vssd1 vccd1 vccd1 _2878_/A sky130_fd_sc_hd__nand4_1
XFILLER_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2703__A1 _4417_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4328_ _4328_/A vssd1 vssd1 vccd1 vccd1 _5327_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input1_A RST_N vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5621__D _5621_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4259_ _4256_/Y _4692_/A _4258_/Y vssd1 vssd1 vccd1 vccd1 _4259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4815__A _4815_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4208__A1 _4147_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4534__B _4550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4253__C _4253_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4550__A _4674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3166__A _3166_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2942__A1 _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input57_A cpu_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__B _4714_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3613__B _3620_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5531__D _5531_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output213_A _3287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4725__A _4725_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3670__A2 _2867_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_CLK clkbuf_1_0_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5798_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5358__CLK _5800_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3630_ _3630_/A _3637_/B _4974_/A vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__and3_1
XANTENNA__4460__A _4891_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3186__A1 input49/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5275__B _5284_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3561_ _4320_/A _5602_/Q _3642_/S vssd1 vssd1 vccd1 vccd1 _4926_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5706__D _5706_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3076__A _4542_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2933__A1 _4423_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5300_ _5300_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5790_/D sky130_fd_sc_hd__nand2_1
X_3492_ _3492_/A vssd1 vssd1 vccd1 vccd1 _3492_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4135__B1 _4134_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5231_ _5231_/A _5266_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__and3_1
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5291__A _5291_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3804__A _4070_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5162_ _5176_/A _5167_/B _5162_/C vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__or3_1
XFILLER_69_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3894__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4113_ _5472_/Q _4074_/X _4112_/X vssd1 vssd1 vccd1 vccd1 _4113_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5441__D _5441_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5093_ _5075_/X _5089_/X _5090_/X _5076_/X _4073_/B vssd1 vssd1 vccd1 vccd1 _5678_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4145_/A _4079_/B _4044_/C vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__and3_1
XFILLER_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3110__A1 _5396_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3661__A2 _4082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5169__C _5184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4946_ _4946_/A vssd1 vssd1 vccd1 vccd1 _5610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4610__A1 _5448_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4073__C _4143_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4610__B2 _4590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2868__B1_N _5694_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4877_ _5268_/A vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4370__A _4378_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3828_ _4692_/A vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__buf_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4801__C _4817_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ _5558_/Q vssd1 vssd1 vccd1 vccd1 _3759_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5616__D _5616_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_3_0_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4126__B1 _4125_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5429_ _5435_/CLK _5429_/D vssd1 vssd1 vccd1 vccd1 _5429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput250 _3391_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput261 _3427_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput272 _3358_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3714__A _3994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput283 _3486_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[10] sky130_fd_sc_hd__buf_2
Xoutput294 _3508_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__2688__B1 _2687_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4529__B _4550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3433__B _3433_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5351__D _5351_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3152__C _4500_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3101__A1 input65/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5500__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4545__A _4674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input111_A ksc_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2860__B1 _2850_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4056__A1_N _3989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5650__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__B1 _2611_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3168__A1 input45/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5526__D _5526_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2915__A1 _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4439__B _4439_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3876__C1 _3875_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3343__B _4761_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output330_A _3621_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__D _5261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3062__C _4460_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5093__A1 _5075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4455__A _4455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2851__B1 _2762_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4174__B _4228_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4800_ _5207_/A vssd1 vssd1 vccd1 vccd1 _4817_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _5798_/CLK _5780_/D vssd1 vssd1 vccd1 vccd1 _5780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2992_ _2994_/A _5428_/Q vssd1 vssd1 vccd1 vccd1 _2993_/A sky130_fd_sc_hd__and2_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4731_ _4731_/A _4731_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__and3_1
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2603__B1 _2916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3800__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4662_ _3756_/X _4667_/C _4266_/Y _4265_/X _4630_/X vssd1 vssd1 vccd1 vccd1 _5483_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3518__B _5653_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3613_ _3613_/A _3620_/B _4959_/C vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__and3_1
XFILLER_50_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5436__D _5436_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _5439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2906__A1 _2829_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3544_ _3558_/A _3547_/B _4911_/A vssd1 vssd1 vccd1 vccd1 _3545_/A sky130_fd_sc_hd__and3_1
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4108__B1 _4107_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5305__C1 _5278_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3475_ _4394_/A _5634_/Q _3654_/S vssd1 vssd1 vccd1 vccd1 _5005_/C sky130_fd_sc_hd__mux2_1
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3534__A _3654_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4659__A1 _5480_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5214_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3867__C1 _3865_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4349__B _4349_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2795__D _2795_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5523__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5145_ _5145_/A _5154_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5146_/A sky130_fd_sc_hd__and3_1
XFILLER_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5076_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4365__A _4365_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3095__A0 _5709_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4027_ _4265_/A vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5673__CLK _5697_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5241__D1 _4429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A vssd1 vssd1 vccd1 vccd1 _5603_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5196__A _5200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3709__A _3709_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2613__A _2622_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5346__D _5346_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3147__C _4498_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3972__A_N _3817_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5311__A2 _5114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input159_A spi_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3086__A0 _4316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4275__A _4287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3610__C _4957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__B1 _2935_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3389__A1 _5506_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4722__B _4731_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4050__A2 _3906_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4441__C _4441_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output280_A _5805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output378_A _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3561__A1 _5602_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5546__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3354__A _3357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2896__C _2909_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _2895_/X _2899_/X _4765_/A vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__o21a_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3073__B _3073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3191_ _5725_/Q input50/X _3223_/S vssd1 vssd1 vccd1 vccd1 _5186_/C sky130_fd_sc_hd__mux2_2
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4266__B1_N _5483_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3864__A2 _3828_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5696__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4185__A _4265_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4813__A1 _5546_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4813__B2 _4804_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2824__B1 _5375_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4913__A _4913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4577__B1 _5807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5763_ _5766_/CLK _5763_/D vssd1 vssd1 vccd1 vccd1 _5763_/Q sky130_fd_sc_hd__dfxtp_1
X_2975_ _5739_/Q input28/X _3233_/S vssd1 vssd1 vccd1 vccd1 _5219_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3529__A _3529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4714_ _4724_/A _4714_/B _4714_/C vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__or3_1
X_5694_ _5694_/CLK _5694_/D vssd1 vssd1 vccd1 vccd1 _5694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4645_ _4645_/A vssd1 vssd1 vccd1 vccd1 _4645_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4576_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4576_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3527_ _3527_/A vssd1 vssd1 vccd1 vccd1 _3527_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3264__A _3453_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3458_ _2924_/X _2927_/X _4990_/C vssd1 vssd1 vccd1 vccd1 _3458_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4079__B _4079_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3389_ _4338_/A _5506_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _4719_/C sky130_fd_sc_hd__mux2_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5128_ _5128_/A _5143_/B _5128_/C vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__or3_1
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4095__A _4110_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5660_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3203__S _3234_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4526__C _4536_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2815__B1 _2932_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4280__A2 _3828_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4823__A _4823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5419__CLK _5695_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4542__B _4542_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4032__A2 _4003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3439__A _3445_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3240__A0 _4292_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5569__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2997__B _5430_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3543__A1 _5597_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3174__A _3174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5296__A1 _5787_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5296__B2 _4104_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3059__A0 _5133_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3113__S _3126_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4271__A2 _3828_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4733__A _4749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4008__C1 _4007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3349__A _3349_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2760_ _5361_/Q vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3068__B _3073_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2691_ _2691_/A vssd1 vssd1 vccd1 vccd1 _2903_/A sky130_fd_sc_hd__clkbuf_4
X_4430_ _5374_/Q _4429_/X _2827_/X _4402_/X vssd1 vssd1 vccd1 vccd1 _5374_/D sky130_fd_sc_hd__a211o_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _5342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5714__D _5714_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3084__A _3174_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3312_ _3314_/A _5547_/Q vssd1 vssd1 vccd1 vccd1 _3313_/A sky130_fd_sc_hd__and2_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4292_ _4299_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__and2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _5124_/C _5314_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__mux2_8
XANTENNA__4908__A _4908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__A2 _3830_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3812__A _4240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3174_/A vssd1 vssd1 vccd1 vccd1 _3219_/S sky130_fd_sc_hd__buf_4
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__C1 _3840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4262__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4362__B _4362_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__A2 _3766_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5711__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5746_ _5767_/CLK _5746_/D vssd1 vssd1 vccd1 vccd1 _5746_/Q sky130_fd_sc_hd__dfxtp_1
X_2958_ _5213_/A _5351_/Q _3229_/S vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__mux2_8
XANTENNA__3773__A1 _3763_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4173__A_N _4075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5677_ _5697_/CLK _5677_/D vssd1 vssd1 vccd1 vccd1 _5677_/Q sky130_fd_sc_hd__dfxtp_1
X_2889_ _2886_/Y _4407_/A _2888_/Y vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__o21ai_4
X_4628_ _4628_/A vssd1 vssd1 vccd1 vccd1 _4667_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5193__B _5202_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4559_ _4559_/A vssd1 vssd1 vccd1 vccd1 _5426_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5624__D _5624_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2610__B _2848_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2733__C1 _2787_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4818__A _4818_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3722__A _4062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4789__B1 _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3461__A0 _4383_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4553__A _4553_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5391__CLK _5435_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3213__A0 _5729_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2567__A2 _2549_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input87_A gpio_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3920__B1_N _5461_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5534__D _5534_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3108__S _3108_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3335__C _4681_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output243_A _5805_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4728__A _4917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3632__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput150 spi_dat_i[15] vssd1 vssd1 vccd1 vccd1 _4043_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput161 spi_dat_i[25] vssd1 vssd1 vccd1 vccd1 _4201_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput172 spi_dat_i[6] vssd1 vssd1 vccd1 vccd1 _3889_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3351__B _3361_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output410_A _3237_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4244__A2 _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5734__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4463__A _4652_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3930_ _3949_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _3930_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3452__B1 _4676_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _4083_/A vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5709__D _5709_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5600_ _5692_/CLK _5600_/D vssd1 vssd1 vccd1 vccd1 _5600_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3204__A0 _4360_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2812_ _4427_/C _4427_/B _4437_/C _4437_/B vssd1 vssd1 vccd1 vccd1 _2816_/C sky130_fd_sc_hd__a22oi_4
XFILLER_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4401__C1 _4379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3792_ _3953_/A _3792_/B _3993_/C _3792_/D vssd1 vssd1 vccd1 vccd1 _3792_/X sky130_fd_sc_hd__and4_2
X_5531_ _5531_/CLK _5531_/D vssd1 vssd1 vccd1 vccd1 _5531_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2558__A2 _5261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2743_ _2698_/A _2640_/X _2742_/Y _2637_/A vssd1 vssd1 vccd1 vccd1 _4437_/B sky130_fd_sc_hd__o211ai_4
XFILLER_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3807__A _3807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2711__A _2711_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ _5482_/CLK _5462_/D vssd1 vssd1 vccd1 vccd1 _5462_/Q sky130_fd_sc_hd__dfxtp_1
X_2674_ _2748_/B _2779_/A _2779_/B _2935_/A vssd1 vssd1 vccd1 vccd1 _2724_/B sky130_fd_sc_hd__and4_1
XANTENNA__3526__B _5657_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4413_ _2591_/Y _2596_/X _4379_/X vssd1 vssd1 vccd1 vccd1 _5364_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__5444__D _5444_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5393_ _5435_/CLK _5393_/D vssd1 vssd1 vccd1 vccd1 _5393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4180__A1 _4147_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4344_ _4344_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__and2_1
XANTENNA__2730__A2 _2645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4638__A _4638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4275_ _4287_/A _4275_/B vssd1 vssd1 vccd1 vccd1 _4275_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3542__A _5058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _3236_/A _4542_/B _4534_/C vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__and3_1
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4357__B _4357_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ _3157_/A vssd1 vssd1 vccd1 vccd1 _3204_/S sky130_fd_sc_hd__buf_2
XFILLER_41_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3691__B1 _2870_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3088_ _3088_/A vssd1 vssd1 vccd1 vccd1 _3088_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__A2 _4229_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4373__A _4373_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4640__C1 _4632_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5619__D _5619_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5729_ _5731_/CLK _5729_/D vssd1 vssd1 vccd1 vccd1 _5729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2621__A _2621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3436__B _3445_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5354__D _5354_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5607__CLK _5692_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2721__A2 _2615_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4548__A _4548_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input141_A ksc_err_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3171__B _3194_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5757__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__A _4283_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__C1 _4630_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4714__C _4714_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A1 _3813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5529__D _5529_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output193_A _4168_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3627__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output360_A _3011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2712__A2 _2549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4458__A _4458_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3362__A _3362_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4060_ _4027_/X _3919_/X _5469_/Q vssd1 vssd1 vccd1 vccd1 _4060_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3081__B _3105_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3011_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4608__D _4614_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3673__B1 _3672_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4870__C1 _4865_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4905__B _4913_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5289__A _5289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3425__A0 _4360_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4962_ _4962_/A vssd1 vssd1 vccd1 vccd1 _5617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3913_ _5776_/Q _3804_/X _3900_/X _3912_/Y vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__3924__B_N _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5439__D _5439_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4893_ _4832_/X _4833_/X _3680_/A _4630_/X vssd1 vssd1 vccd1 vccd1 _5589_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4921__A _4921_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3844_ _4091_/A vssd1 vssd1 vccd1 vccd1 _5268_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3775_ _4628_/A _3756_/X _5099_/A _3774_/Y vssd1 vssd1 vccd1 vccd1 _3775_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3537__A _3537_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2936__C1 _2935_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5514_ _5694_/CLK _5514_/D vssd1 vssd1 vccd1 vccd1 _5514_/Q sky130_fd_sc_hd__dfxtp_1
X_2726_ _2726_/A vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__buf_2
X_5445_ _5531_/CLK _5445_/D vssd1 vssd1 vccd1 vccd1 _5445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput410 _3237_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[31] sky130_fd_sc_hd__buf_2
X_2657_ _2695_/C _2695_/D _2695_/B _5759_/Q vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__a31o_2
Xoutput421 _3253_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_47_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5376_ _5765_/CLK _5376_/D vssd1 vssd1 vccd1 vccd1 _5376_/Q sky130_fd_sc_hd__dfxtp_2
X_2588_ _2572_/Y _2574_/X _2587_/Y vssd1 vssd1 vccd1 vccd1 _4411_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__2703__A2 _4417_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4327_ _4344_/A _4327_/B vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__and2_1
XANTENNA__4368__A _4368_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4258_ _3763_/A _3766_/A _3768_/A _4257_/X _4117_/A vssd1 vssd1 vccd1 vccd1 _4258_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_68_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3209_ _4362_/B _5413_/Q _3209_/S vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__mux2_1
X_4189_ _3860_/X _3861_/X _4189_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _4189_/X sky130_fd_sc_hd__and4bb_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4208__A2 _3722_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5199__A _5199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__A _2616_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4613__C1 _4598_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4534__C _4534_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5349__D _5349_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4253__D _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4831__A _4831_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4550__B _4550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2942__A2 _2927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__C _4709_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3613__C _4959_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3655__B1 _4905_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4852__C1 _4840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output206_A _3882_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3121__S _3132_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4080__B1 _4079_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__A _4741_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4460__B _4473_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3357__A _3357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3560_ _5058_/A vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4239__A1_N _3806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2933__A2 _4423_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3491_ _3493_/A _5641_/Q vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__and2_1
XFILLER_66_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5230_ _2614_/Y _5227_/A _2618_/Y vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4135__A1 _4059_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5291__B _5297_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _5161_/A vssd1 vssd1 vccd1 vccd1 _5714_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4188__A _5581_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5722__D _5722_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3092__A _3092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3894__B1 _3892_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4112_ _4145_/A _4228_/B _4112_/C vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__and3_2
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _5081_/X _5078_/X _5087_/X _5084_/X _4058_/B vssd1 vssd1 vccd1 vccd1 _5677_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4043_ _3817_/X _3818_/X _4043_/C _4043_/D vssd1 vssd1 vccd1 vccd1 _4044_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__4916__A _4916_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3661__A3 _4083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4945_ _4963_/A _4963_/B _4945_/C vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__or3_1
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4610__A2 _4573_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4073__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4651__A _4651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4876_ _5089_/A vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5452__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3827_ _5560_/Q vssd1 vssd1 vccd1 vccd1 _3827_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3267__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3758_ _3758_/A vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2616_/X _2617_/X _5765_/Q vssd1 vssd1 vccd1 vccd1 _2709_/Y sky130_fd_sc_hd__o21bai_4
X_3689_ _4153_/A vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__buf_2
X_5428_ _5435_/CLK _5428_/D vssd1 vssd1 vccd1 vccd1 _5428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4126__B2 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput240 _3276_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[7] sky130_fd_sc_hd__buf_2
Xoutput251 _3394_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput262 _3430_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput273 _3362_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput284 _3488_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2688__A1 _5758_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5359_ _5800_/CLK _5359_/D vssd1 vssd1 vccd1 vccd1 _5359_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4098__A _4098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput295 _3510_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[21] sky130_fd_sc_hd__buf_2
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5632__D _5632_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4529__C _4529_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3433__C _4749_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4826__A _4826_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3730__A _3980_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4834__C1 _4630_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4545__B _4550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2860__A1 _2751_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input104_A gpio_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4561__A _4561_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2612__A1 _2605_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4257__A_N _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3177__A _3183_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2915__A2 _2899_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3905__A _5564_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3624__B _3637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5542__D _5542_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3116__S _3151_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3876__B1 _5099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4439__C _4439_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3343__C _4686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5325__CLK _5766_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2955__S _3228_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4736__A _4947_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output323_A _3599_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3640__A _3646_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5093__A2 _5089_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2851__A1 _2760_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5475__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4174__C _4174_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ _3029_/A vssd1 vssd1 vccd1 vccd1 _2994_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__B1 _4041_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4471__A _4471_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4730_ _4730_/A vssd1 vssd1 vccd1 vccd1 _5510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2603__A1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__B1 _3798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4661_ _5482_/Q _4652_/X _4254_/X _4621_/A vssd1 vssd1 vccd1 vccd1 _5482_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5717__D _5717_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3087__A _3092_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3612_ _4351_/A _5616_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _4959_/C sky130_fd_sc_hd__mux2_1
XFILLER_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4592_ _4592_/A _5439_/Q _4604_/C _4596_/D vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__and4_1
XFILLER_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2906__A2 _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3543_ _4308_/B _5597_/Q _3564_/S vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3815__A _4489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5305__B1 _4214_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4108__B2 _3934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3474_ _3469_/X _3470_/X _5003_/A vssd1 vssd1 vccd1 vccd1 _3474_/X sky130_fd_sc_hd__o21a_1
XFILLER_100_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4659__A2 _4652_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5213_ _5213_/A _5225_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__and3_1
XANTENNA__5452__D _5452_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3867__B1 _3856_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5144_ _5144_/A vssd1 vssd1 vccd1 vccd1 _5707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3619__A0 _4355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4816__C1 _4805_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3550__A _4988_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4026_ _4127_/A _4026_/B _4159_/C _4026_/D vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__and4_2
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3095__A1 input64/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4084__C _4084_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5241__C1 _5228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4381__A _4381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4928_ _4928_/A _4940_/B _4940_/C vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__and3_1
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5196__B _5215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5627__D _5627_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4859_ _5081_/A vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3725__A _4781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5348__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5362__D _5362_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5311__A3 _5069_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4556__A _4556_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3460__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5498__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3086__A1 _5392_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4275__B _4275_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__A1 _2829_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4035__B1 _4026_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4291__A _4441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4722__C _4741_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5537__D _5537_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2671__A_N input20/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3797__A_N _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output273_A _3362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3635__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2896__D _2929_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3354__B _3361_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3073__C _4469_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3190_/A vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4466__A _4466_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3370__A _3370_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4274__B1 _4273_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4185__B _4265_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4813__A2 _4803_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2824__A1 _2806_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4913__B _4913_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5297__A _5297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4577__A1 _5432_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5762_ _5767_/CLK _5762_/D vssd1 vssd1 vccd1 vccd1 _5762_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4577__B2 _4564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2974_ _4295_/B vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2588__B1 _2587_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4713_ _4713_/A vssd1 vssd1 vccd1 vccd1 _5503_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5447__D _5447_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5693_ _5694_/CLK _5693_/D vssd1 vssd1 vccd1 vccd1 _5693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4644_ _4651_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _5467_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4575_ _5204_/A vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__buf_4
XANTENNA__3545__A _3545_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3526_ _3526_/A _5657_/Q vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__and2_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3457_ _4381_/A _5628_/Q _3645_/S vssd1 vssd1 vccd1 vccd1 _4990_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4079__C _4079_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5640__CLK _5659_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3388_ _3388_/A vssd1 vssd1 vccd1 vccd1 _3388_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5127_ _5127_/A vssd1 vssd1 vccd1 vccd1 _5700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4376__A _5212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3280__A _3280_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5058_ _5058_/A _5058_/B _5235_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__and3_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _5781_/Q _3915_/X _3993_/X _4008_/Y vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__o22ai_4
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5790__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2815__A1 _2565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4017__B1 _4016_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2624__A _2686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4542__C _5266_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5000__A _5000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3439__B _3445_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3240__A1 _5383_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5357__D _5357_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3455__A _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input171_A spi_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5296__A2 _5289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A cpu_adr_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3190__A _3190_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3059__A1 _5318_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4008__B1 _4006_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4733__B _4739_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output390_A _3135_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5513__CLK _5555_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3068__C _4464_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2690_ _5379_/Q vssd1 vssd1 vccd1 vccd1 _2690_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2990__B1 _4561_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3365__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4192__C1 _4191_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4360_ _4360_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__or2_1
XANTENNA__5663__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3311_ _3311_/A vssd1 vssd1 vccd1 vccd1 _3311_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2742__B1 _5764_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4291_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__clkbuf_4
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _5699_/Q input68/X _3250_/S vssd1 vssd1 vccd1 vccd1 _5124_/C sky130_fd_sc_hd__mux2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3812__B _3812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3173_ _5722_/Q input47/X _3186_/S vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4196__A _4196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5730__D _5730_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4247__B1 _4246_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4924__A _4924_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5745_ _5767_/CLK _5745_/D vssd1 vssd1 vccd1 vccd1 _5745_/Q sky130_fd_sc_hd__dfxtp_1
X_2957_ _3174_/A vssd1 vssd1 vccd1 vccd1 _3229_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3773__A2 _3766_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2888_ _2631_/Y _2724_/Y _5419_/Q vssd1 vssd1 vccd1 vccd1 _2888_/Y sky130_fd_sc_hd__o21ai_1
X_5676_ _5694_/CLK _5676_/D vssd1 vssd1 vccd1 vccd1 _5676_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2981__A0 _4392_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4627_ _5456_/Q _4623_/X _3821_/X _4660_/A vssd1 vssd1 vccd1 vccd1 _5456_/D sky130_fd_sc_hd__a211o_1
XFILLER_85_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5193__C _5208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4558_ _4674_/A _4558_/B _4558_/C vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__or3_1
XANTENNA__2610__C _2848_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2733__B1 _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3509_ _3515_/A _5649_/Q vssd1 vssd1 vccd1 vccd1 _3510_/A sky130_fd_sc_hd__and2_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__buf_2
XFILLER_46_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__D _5640_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3214__S _3234_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4789__A1 _5534_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4789__B2 _4782_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3461__A1 _5629_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5536__CLK _5538_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3749__C1 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3213__A1 input54/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5686__CLK _5690_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2972__B1 _4552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3185__A _3212_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3835__A_N _3832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput140 ksc_dat_i[9] vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5550__D _5550_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output236_A _3266_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput151 spi_dat_i[16] vssd1 vssd1 vccd1 vccd1 _4061_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput162 spi_dat_i[26] vssd1 vssd1 vccd1 vccd1 _4216_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput173 spi_dat_i[7] vssd1 vssd1 vccd1 vccd1 _3902_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3351__C _4690_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4229__B1 _4228_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2963__S _3233_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output403_A _3206_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4744__A _4749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3452__A1 _3281_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3860_ _4082_/A vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2811_ _2809_/X _2676_/X _2690_/Y vssd1 vssd1 vccd1 vccd1 _4437_/C sky130_fd_sc_hd__o21ai_4
XANTENNA__3204__A1 _5412_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ _4171_/A vssd1 vssd1 vccd1 vccd1 _3993_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4401__B1 _2619_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5530_ _5538_/CLK _5530_/D vssd1 vssd1 vccd1 vccd1 _5530_/Q sky130_fd_sc_hd__dfxtp_1
X_2742_ _2616_/X _2617_/X _5764_/Q vssd1 vssd1 vccd1 vccd1 _2742_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2963__A0 _5737_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _5741_/CLK _5461_/D vssd1 vssd1 vccd1 vccd1 _5461_/Q sky130_fd_sc_hd__dfxtp_1
X_2673_ _5761_/Q _2577_/X _2671_/Y _2704_/A _2806_/A vssd1 vssd1 vccd1 vccd1 _2935_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5725__D _5725_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4412_ _4412_/A vssd1 vssd1 vccd1 vccd1 _5363_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4165__C1 _4835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5392_ _5731_/CLK _5392_/D vssd1 vssd1 vccd1 vccd1 _5392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4343_ _4343_/A vssd1 vssd1 vccd1 vccd1 _5334_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3912__C1 _3840_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4180__A2 _4046_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__A _5005_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3823__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5409__CLK _5446_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4274_ _5799_/Q _3690_/X _4273_/Y vssd1 vssd1 vccd1 vccd1 _4275_/B sky130_fd_sc_hd__o21ai_4
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4638__B _4638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3225_ _4368_/A _5416_/Q _3235_/S vssd1 vssd1 vccd1 vccd1 _4534_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5460__D _5460_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3140__A0 _4335_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3156_ _5172_/C _5334_/Q _3192_/S vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__mux2_8
XANTENNA__3691__A1 _5694_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5559__CLK _5802_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4654__A _4660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3087_ _3092_/A _3105_/B _4473_/C vssd1 vssd1 vccd1 vccd1 _3088_/A sky130_fd_sc_hd__and3_1
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4373__B _4381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4640__B1 _3973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _3989_/X sky130_fd_sc_hd__buf_2
XANTENNA__2902__A _2902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5728_ _5731_/CLK _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5659_ _5659_/CLK _5659_/D vssd1 vssd1 vccd1 vccd1 _5659_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5635__D _5635_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3209__S _3209_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3436__C _4751_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2706__B1 _2705_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4829__A _4829_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4548__B _4556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5370__D _5370_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3131__A0 _5715_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3171__C _4510_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A ksc_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4564__A _4590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__B _4283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__B1 _3853_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3985__A2 _3974_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__C1 _2574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3198__A0 _5189_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__A _4117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2945__A0 _5735_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3627__B _3637_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5545__D _5545_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output186_A _4069_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2958__S _3229_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output353_A _2952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4739__A _4749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3643__A _3646_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__A_N _3860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4458__B _4475_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5701__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4177__C _4177_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3122__A0 _4329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3010_ _3016_/A _5436_/Q vssd1 vssd1 vccd1 vccd1 _3011_/A sky130_fd_sc_hd__and2_1
XANTENNA__3081__C _4471_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3673__A1 _4139_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4870__B1 _4856_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4474__A _4474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4905__C _4905_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _4961_/A _4965_/B _4965_/C vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__and3_1
XANTENNA__3425__A1 _5516_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3912_ _3813_/X _3904_/Y _3911_/Y _3840_/X vssd1 vssd1 vccd1 vccd1 _3912_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4892_ _4889_/X _4890_/X _4280_/Y _4891_/X vssd1 vssd1 vccd1 vccd1 _5588_/D sky130_fd_sc_hd__a211o_1
XFILLER_60_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3843_ _3869_/A _5277_/A vssd1 vssd1 vccd1 vccd1 _3843_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3818__A _4076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3774_ _3759_/Y _4743_/A _3773_/Y vssd1 vssd1 vccd1 vccd1 _3774_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2936__B1 _2821_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5513_ _5555_/CLK _5513_/D vssd1 vssd1 vccd1 vccd1 _5513_/Q sky130_fd_sc_hd__dfxtp_1
X_2725_ _2631_/Y _2724_/Y _2561_/Y vssd1 vssd1 vccd1 vccd1 _2726_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__5455__D _5455_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5444_ _5446_/CLK _5444_/D vssd1 vssd1 vccd1 vccd1 _5444_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput400 _3190_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[22] sky130_fd_sc_hd__buf_2
X_2656_ _2780_/A _2782_/A _2780_/C _2782_/B vssd1 vssd1 vccd1 vccd1 _2724_/A sky130_fd_sc_hd__and4_1
Xoutput411 _3074_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput422 _5807_/X vssd1 vssd1 vccd1 vccd1 spi_stb_o sky130_fd_sc_hd__buf_2
XFILLER_47_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2587_ _5748_/Q _2577_/X _2585_/Y _2696_/A vssd1 vssd1 vccd1 vccd1 _2587_/Y sky130_fd_sc_hd__o211ai_1
X_5375_ _5741_/CLK _5375_/D vssd1 vssd1 vccd1 vccd1 _5375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4649__A _4651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3553__A _3553_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4326_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4368__B _4381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5381__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _3999_/A _4000_/A _4257_/C _4257_/D vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__and4bb_2
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3113__A0 _5712_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3208_ _5193_/A _5343_/Q _3219_/S vssd1 vssd1 vccd1 vccd1 _4362_/B sky130_fd_sc_hd__mux2_8
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4188_ _5581_/Q vssd1 vssd1 vccd1 vccd1 _4188_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3139_ _5165_/A _5331_/Q _3162_/S vssd1 vssd1 vccd1 vccd1 _4335_/B sky130_fd_sc_hd__mux2_8
XANTENNA__4384__A _4384_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4613__B1 _3062_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3728__A _4083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2632__A _5372_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4550__C _4550_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5365__D _5365_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4559__A _4559_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5724__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3104__A0 _4322_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3655__A1 _3482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4852__B1 _3910_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4294__A input1/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__A1 _5470_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4741__B _4756_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__A _3638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2542__A _5768_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4460__C _4460_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3357__B _3361_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2918__B1 _5660_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _3490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4135__A2 _4651_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4469__A _4487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3373__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5160_ _5160_/A _5178_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__and3_1
XFILLER_97_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3894__A1 _3720_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3092__B _3105_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3894__B2 _3893_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4111_ _4075_/X _4076_/X _4111_/C _4201_/D vssd1 vssd1 vccd1 vccd1 _4112_/C sky130_fd_sc_hd__and4bb_1
X_5091_ _5075_/X _5089_/X _5090_/X _5076_/X _4041_/B vssd1 vssd1 vccd1 vccd1 _5676_/D
+ sky130_fd_sc_hd__a311o_1
X_4042_ _4059_/A vssd1 vssd1 vccd1 vccd1 _4042_/X sky130_fd_sc_hd__buf_2
XANTENNA__4096__B1_N _5471_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4932__A _4932_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4944_ _5005_/B vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4651__B _4651_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4875_ _5081_/A vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3548__A _3548_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3826_ _4005_/A vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__buf_2
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5747__CLK _5767_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3757_ _3757_/A vssd1 vssd1 vccd1 vccd1 _3758_/A sky130_fd_sc_hd__buf_2
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2708_ _2708_/A vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__clkbuf_4
X_3688_ _3742_/A vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_12_CLK_A clkbuf_1_1_1_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput230 _3322_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[27] sky130_fd_sc_hd__buf_2
X_5427_ _5435_/CLK _5427_/D vssd1 vssd1 vccd1 vccd1 _5427_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4379__A _4431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2639_ _2639_/A vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__inv_2
Xoutput241 _3280_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[8] sky130_fd_sc_hd__buf_2
XANTENNA__3283__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3334__A0 _4304_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput252 _3398_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput263 _3434_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput274 _3366_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_82_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput285 _3490_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[12] sky130_fd_sc_hd__buf_2
X_5358_ _5800_/CLK _5358_/D vssd1 vssd1 vccd1 vccd1 _5358_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2688__A2 _2683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput296 _3512_/X vssd1 vssd1 vccd1 vccd1 ksc_adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _5319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5289_ _5289_/A vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4834__B1 _4832_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5003__A _5003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4545__C _4545_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2860__A2 _2574_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4842__A _4971_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4561__B _4681_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__A2 _2606_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3177__B _3194_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3573__A0 _4327_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3888__B1_N _5459_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input62_A cpu_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3624__C _4965_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3876__A1 _4628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3640__B _4988_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5093__A3 _5090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output316_A _3575_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3132__S _3132_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2851__A2 _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2971__S _3240_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4752__A _4752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4053__A1 _5784_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2990_ _2973_/X _2974_/X _4561_/A vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__o21a_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__B1 _5242_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__B2 _4052_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4201__A_N _4075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__B _4475_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2603__A2 _2596_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3800__A1 _3720_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3800__B2 _3799_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4660_ _4660_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _5481_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3087__B _3105_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4591_ _5438_/Q _4589_/X _4584_/X _4590_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _5438_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3564__A0 _4322_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3542_ _5058_/A vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5305__A1 _5795_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3473_ _4392_/B _5633_/Q _3652_/S vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5305__B2 _4221_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4199__A _4199_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5733__D _5733_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5212_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5231_/C sky130_fd_sc_hd__buf_2
XFILLER_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3867__A1 _5072_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5143_ _5152_/A _5143_/B _5143_/C vssd1 vssd1 vccd1 vccd1 _5144_/A sky130_fd_sc_hd__or3_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4927__A _4927_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3831__A _3979_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5074_ _4889_/X _5060_/X _5066_/X _5061_/X _3886_/B vssd1 vssd1 vccd1 vccd1 _5667_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3619__A1 _5618_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4816__B1 _4798_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4025_ _4171_/A vssd1 vssd1 vccd1 vccd1 _4159_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__2827__C1 _2574_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4084__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5241__B1 _2595_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _5602_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4381__B _4381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3278__A _3316_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5196__C _5196_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4858_ _3960_/X _3962_/X _4856_/X _4857_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _5567_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3809_ _3806_/X _5664_/Q _3807_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _3812_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789_ _5534_/Q _4780_/X _5805_/A _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _5534_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2910__A _2910_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3937__B_N _3818_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5643__D _5643_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4837__A _4837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4556__B _4556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__A2 _2565_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4572__A _4595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4035__A1 _5783_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4035__B2 _4034_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3546__A0 _4310_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3916__A _3916_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5553__D _5553_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output266_A _3344_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3127__S _3162_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3354__C _4694_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2966__S _3235_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4747__A _4747_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5442__CLK _5531_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4274__A1 _5799_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4185__C _4265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2824__A2 _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5592__CLK _5635_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4482__A _4482_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4913__C _4913_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5297__B _5297_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4577__A2 _4563_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5761_ _5765_/CLK _5761_/D vssd1 vssd1 vccd1 vccd1 _5761_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _3042_/A vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5728__D _5728_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2588__A1 _2572_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4712_ _4712_/A _4731_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__and3_1
XANTENNA__3785__B1 _5289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5692_ _5692_/CLK _5692_/D vssd1 vssd1 vccd1 vccd1 _5692_/Q sky130_fd_sc_hd__dfxtp_1
X_4643_ _5466_/Q _4639_/X _4018_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _5466_/D sky130_fd_sc_hd__a211o_1
XFILLER_50_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3826__A _4005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4574_ _4574_/A vssd1 vssd1 vccd1 vccd1 _5431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3525_ _3525_/A vssd1 vssd1 vccd1 vccd1 _3525_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3891__A_N _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5463__D _5463_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3456_ _4289_/D vssd1 vssd1 vccd1 vccd1 _3645_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3387_ _3393_/A _3397_/B _4716_/A vssd1 vssd1 vccd1 vccd1 _3388_/A sky130_fd_sc_hd__and3_1
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5126_ _5126_/A _5130_/B _5236_/A vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__and3_1
XFILLER_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5057_ _5057_/A vssd1 vssd1 vccd1 vccd1 _5659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4008_ _3887_/X _4642_/B _4006_/Y _4007_/X vssd1 vssd1 vccd1 vccd1 _4008_/Y sky130_fd_sc_hd__o211ai_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2815__A2 _2677_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4392__A _4396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4017__A1 _4011_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5638__D _5638_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3776__B1 _3775_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3439__C _4754_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5315__CLK _5765_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3736__A _3736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2640__A _2640_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5373__D _5373_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5465__CLK _5482_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input164_A spi_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4567__A _4567_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3902__C _3902_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input25_A cpu_adr_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4008__A1 _3887_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4733__C _4733_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5548__D _5548_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output383_A _2993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3646__A _3646_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2990__A1 _2973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3365__B _3380_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4192__B1 _3826_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2742__A1 _2616_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3310_ _3314_/A _5546_/Q vssd1 vssd1 vccd1 vccd1 _3311_/A sky130_fd_sc_hd__and2_1
X_4290_ _4378_/A vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__clkbuf_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3241_ _2973_/X _2974_/X _4445_/A vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__o21a_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4477__A _4558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3381__A _3381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _3172_/A vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3812__C _4240_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A1 _3813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4924__B _4940_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5458__D _5458_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5338__CLK _5737_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4940__A _4940_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5744_ _5766_/CLK _5744_/D vssd1 vssd1 vccd1 vccd1 _5744_/Q sky130_fd_sc_hd__dfxtp_1
X_2956_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3174_/A sky130_fd_sc_hd__buf_2
XFILLER_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5675_ _5697_/CLK _5675_/D vssd1 vssd1 vccd1 vccd1 _5675_/Q sky130_fd_sc_hd__dfxtp_1
X_2887_ _2909_/A _2925_/A _2887_/C _2925_/B vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__nand4_4
XANTENNA__3556__A _3556_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2981__A1 _5425_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5488__CLK _5586_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4626_ _4638_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _5455_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3657__B1_N _2845_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4557_ _4557_/A vssd1 vssd1 vccd1 vccd1 _5425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2610__D _2848_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2733__A1 _4415_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3508_ _3508_/A vssd1 vssd1 vccd1 vccd1 _3508_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4488_ _4488_/A vssd1 vssd1 vccd1 vccd1 _5398_/D sky130_fd_sc_hd__clkbuf_1
X_3439_ _3445_/A _3445_/B _4754_/C vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__and3_1
XANTENNA__4387__A _4387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3291__A _3291_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5099_/X _5094_/X _5066_/A _5102_/X _4240_/B vssd1 vssd1 vccd1 vccd1 _5689_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4789__A2 _4780_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2635__A _2686_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__S _3230_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__5011__A _5034_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5368__D _5368_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3749__B1 _5058_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3466__A _3654_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2972__A1 _2876_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3921__B1 _3920_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4297__A _4297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput130 ksc_dat_i[29] vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 ksc_err_i vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput152 spi_dat_i[17] vssd1 vssd1 vccd1 vccd1 _4078_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput163 spi_dat_i[27] vssd1 vssd1 vccd1 vccd1 _4227_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput174 spi_dat_i[8] vssd1 vssd1 vccd1 vccd1 _3921_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__4229__A1 _5480_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output229_A _3320_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4744__B _4763_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2545__A _2640_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3140__S _3151_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3452__A2 _2899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4760__A _4947_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2810_ _2809_/X _2750_/X _2682_/Y vssd1 vssd1 vccd1 vccd1 _4427_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__4401__A1 _5359_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5630__CLK _5694_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2741_ _2741_/A _2741_/B vssd1 vssd1 vccd1 vccd1 _2877_/A sky130_fd_sc_hd__nor2_4
XANTENNA__3376__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2963__A1 input24/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_CLK clkbuf_1_1_1_CLK/X vssd1 vssd1 vccd1 vccd1 _5692_/CLK sky130_fd_sc_hd__clkbuf_16
X_5460_ _5482_/CLK _5460_/D vssd1 vssd1 vccd1 vccd1 _5460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2672_ _2672_/A vssd1 vssd1 vccd1 vccd1 _2806_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4411_ _4573_/D _5102_/A _4411_/C vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__and3_1
XANTENNA__4165__B1 _4163_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_5391_ _5435_/CLK _5391_/D vssd1 vssd1 vccd1 vccd1 _5391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5780__CLK _5798_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3912__B1 _3911_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4342_ _4342_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__or2_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__5741__D _5741_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4273_ _5111_/A _3848_/X _4267_/Y _4272_/Y _3866_/X vssd1 vssd1 vccd1 vccd1 _4273_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_84_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4000__A _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3224_ _5200_/C _5346_/Q _3234_/S vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__mux2_8
.ends

