* NGSPICE file created from mkQF100Fabric.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__fakediode_2 abstract view
.subckt sky130_ef_sc_hd__fakediode_2 DIODE VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt mkQF100Fabric CLK RST_N cpu_ack_o cpu_adr_i[0] cpu_adr_i[10] cpu_adr_i[11]
+ cpu_adr_i[12] cpu_adr_i[13] cpu_adr_i[14] cpu_adr_i[15] cpu_adr_i[16] cpu_adr_i[17]
+ cpu_adr_i[18] cpu_adr_i[19] cpu_adr_i[1] cpu_adr_i[20] cpu_adr_i[21] cpu_adr_i[22]
+ cpu_adr_i[23] cpu_adr_i[24] cpu_adr_i[25] cpu_adr_i[26] cpu_adr_i[27] cpu_adr_i[28]
+ cpu_adr_i[29] cpu_adr_i[2] cpu_adr_i[30] cpu_adr_i[31] cpu_adr_i[3] cpu_adr_i[4]
+ cpu_adr_i[5] cpu_adr_i[6] cpu_adr_i[7] cpu_adr_i[8] cpu_adr_i[9] cpu_cyc_i cpu_dat_i[0]
+ cpu_dat_i[10] cpu_dat_i[11] cpu_dat_i[12] cpu_dat_i[13] cpu_dat_i[14] cpu_dat_i[15]
+ cpu_dat_i[16] cpu_dat_i[17] cpu_dat_i[18] cpu_dat_i[19] cpu_dat_i[1] cpu_dat_i[20]
+ cpu_dat_i[21] cpu_dat_i[22] cpu_dat_i[23] cpu_dat_i[24] cpu_dat_i[25] cpu_dat_i[26]
+ cpu_dat_i[27] cpu_dat_i[28] cpu_dat_i[29] cpu_dat_i[2] cpu_dat_i[30] cpu_dat_i[31]
+ cpu_dat_i[3] cpu_dat_i[4] cpu_dat_i[5] cpu_dat_i[6] cpu_dat_i[7] cpu_dat_i[8] cpu_dat_i[9]
+ cpu_dat_o[0] cpu_dat_o[10] cpu_dat_o[11] cpu_dat_o[12] cpu_dat_o[13] cpu_dat_o[14]
+ cpu_dat_o[15] cpu_dat_o[16] cpu_dat_o[17] cpu_dat_o[18] cpu_dat_o[19] cpu_dat_o[1]
+ cpu_dat_o[20] cpu_dat_o[21] cpu_dat_o[22] cpu_dat_o[23] cpu_dat_o[24] cpu_dat_o[25]
+ cpu_dat_o[26] cpu_dat_o[27] cpu_dat_o[28] cpu_dat_o[29] cpu_dat_o[2] cpu_dat_o[30]
+ cpu_dat_o[31] cpu_dat_o[3] cpu_dat_o[4] cpu_dat_o[5] cpu_dat_o[6] cpu_dat_o[7] cpu_dat_o[8]
+ cpu_dat_o[9] cpu_err_o cpu_rty_o cpu_sel_i[0] cpu_sel_i[1] cpu_sel_i[2] cpu_sel_i[3]
+ cpu_stb_i cpu_we_i gpio_ack_i gpio_adr_o[0] gpio_adr_o[10] gpio_adr_o[11] gpio_adr_o[12]
+ gpio_adr_o[13] gpio_adr_o[14] gpio_adr_o[15] gpio_adr_o[16] gpio_adr_o[17] gpio_adr_o[18]
+ gpio_adr_o[19] gpio_adr_o[1] gpio_adr_o[20] gpio_adr_o[21] gpio_adr_o[22] gpio_adr_o[23]
+ gpio_adr_o[24] gpio_adr_o[25] gpio_adr_o[26] gpio_adr_o[27] gpio_adr_o[28] gpio_adr_o[29]
+ gpio_adr_o[2] gpio_adr_o[30] gpio_adr_o[31] gpio_adr_o[3] gpio_adr_o[4] gpio_adr_o[5]
+ gpio_adr_o[6] gpio_adr_o[7] gpio_adr_o[8] gpio_adr_o[9] gpio_cyc_o gpio_dat_i[0]
+ gpio_dat_i[10] gpio_dat_i[11] gpio_dat_i[12] gpio_dat_i[13] gpio_dat_i[14] gpio_dat_i[15]
+ gpio_dat_i[16] gpio_dat_i[17] gpio_dat_i[18] gpio_dat_i[19] gpio_dat_i[1] gpio_dat_i[20]
+ gpio_dat_i[21] gpio_dat_i[22] gpio_dat_i[23] gpio_dat_i[24] gpio_dat_i[25] gpio_dat_i[26]
+ gpio_dat_i[27] gpio_dat_i[28] gpio_dat_i[29] gpio_dat_i[2] gpio_dat_i[30] gpio_dat_i[31]
+ gpio_dat_i[3] gpio_dat_i[4] gpio_dat_i[5] gpio_dat_i[6] gpio_dat_i[7] gpio_dat_i[8]
+ gpio_dat_i[9] gpio_dat_o[0] gpio_dat_o[10] gpio_dat_o[11] gpio_dat_o[12] gpio_dat_o[13]
+ gpio_dat_o[14] gpio_dat_o[15] gpio_dat_o[16] gpio_dat_o[17] gpio_dat_o[18] gpio_dat_o[19]
+ gpio_dat_o[1] gpio_dat_o[20] gpio_dat_o[21] gpio_dat_o[22] gpio_dat_o[23] gpio_dat_o[24]
+ gpio_dat_o[25] gpio_dat_o[26] gpio_dat_o[27] gpio_dat_o[28] gpio_dat_o[29] gpio_dat_o[2]
+ gpio_dat_o[30] gpio_dat_o[31] gpio_dat_o[3] gpio_dat_o[4] gpio_dat_o[5] gpio_dat_o[6]
+ gpio_dat_o[7] gpio_dat_o[8] gpio_dat_o[9] gpio_err_i gpio_rty_i gpio_sel_o[0] gpio_sel_o[1]
+ gpio_sel_o[2] gpio_sel_o[3] gpio_stb_o gpio_we_o spi_ack_i spi_adr_o[0] spi_adr_o[10]
+ spi_adr_o[11] spi_adr_o[12] spi_adr_o[13] spi_adr_o[14] spi_adr_o[15] spi_adr_o[16]
+ spi_adr_o[17] spi_adr_o[18] spi_adr_o[19] spi_adr_o[1] spi_adr_o[20] spi_adr_o[21]
+ spi_adr_o[22] spi_adr_o[23] spi_adr_o[24] spi_adr_o[25] spi_adr_o[26] spi_adr_o[27]
+ spi_adr_o[28] spi_adr_o[29] spi_adr_o[2] spi_adr_o[30] spi_adr_o[31] spi_adr_o[3]
+ spi_adr_o[4] spi_adr_o[5] spi_adr_o[6] spi_adr_o[7] spi_adr_o[8] spi_adr_o[9] spi_cyc_o
+ spi_dat_i[0] spi_dat_i[10] spi_dat_i[11] spi_dat_i[12] spi_dat_i[13] spi_dat_i[14]
+ spi_dat_i[15] spi_dat_i[16] spi_dat_i[17] spi_dat_i[18] spi_dat_i[19] spi_dat_i[1]
+ spi_dat_i[20] spi_dat_i[21] spi_dat_i[22] spi_dat_i[23] spi_dat_i[24] spi_dat_i[25]
+ spi_dat_i[26] spi_dat_i[27] spi_dat_i[28] spi_dat_i[29] spi_dat_i[2] spi_dat_i[30]
+ spi_dat_i[31] spi_dat_i[3] spi_dat_i[4] spi_dat_i[5] spi_dat_i[6] spi_dat_i[7] spi_dat_i[8]
+ spi_dat_i[9] spi_dat_o[0] spi_dat_o[10] spi_dat_o[11] spi_dat_o[12] spi_dat_o[13]
+ spi_dat_o[14] spi_dat_o[15] spi_dat_o[16] spi_dat_o[17] spi_dat_o[18] spi_dat_o[19]
+ spi_dat_o[1] spi_dat_o[20] spi_dat_o[21] spi_dat_o[22] spi_dat_o[23] spi_dat_o[24]
+ spi_dat_o[25] spi_dat_o[26] spi_dat_o[27] spi_dat_o[28] spi_dat_o[29] spi_dat_o[2]
+ spi_dat_o[30] spi_dat_o[31] spi_dat_o[3] spi_dat_o[4] spi_dat_o[5] spi_dat_o[6]
+ spi_dat_o[7] spi_dat_o[8] spi_dat_o[9] spi_err_i spi_rty_i spi_sel_o[0] spi_sel_o[1]
+ spi_sel_o[2] spi_sel_o[3] spi_stb_o spi_we_o vccd1 vssd1
XANTENNA__2479__B1 _2473_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4357__D _4357_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3691__A2 _3351_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _3174_/B _4182_/Q _3206_/A vssd1 vssd1 vccd1 vccd1 _3572_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2158__C _2158_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3086_ _3099_/A _3089_/B _3609_/A vssd1 vssd1 vccd1 vccd1 _3087_/A sky130_fd_sc_hd__and3_1
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2106_ _2106_/A vssd1 vssd1 vccd1 vccd1 _2129_/B sky130_fd_sc_hd__buf_2
XANTENNA__2455__A _4261_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3979__B1 _2489_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2037_ _2037_/A vssd1 vssd1 vccd1 vccd1 _2038_/A sky130_fd_sc_hd__clkinv_2
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4092__D _4092_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3988_ _3952_/X _3955_/X _2569_/Y vssd1 vssd1 vccd1 vccd1 _4379_/D sky130_fd_sc_hd__o21bai_1
X_2939_ _2939_/A vssd1 vssd1 vccd1 vccd1 _2939_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2403__B1 _2239_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3717__C _3721_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3286__A _3328_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2954__A1 _4009_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4108__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4258__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3131__A1 _4210_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4267__D _4267_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input127_A spi_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2365__A _4257_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__B1 _4002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2084__B _2084_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input92_A gpio_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2812__B _2812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3196__A _3196_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2945__A1 input67/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output179_A _2996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2173__A2 _2001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4177__D _4177_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4389_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2881__A0 _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2275__A _2412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2633__B1 _2469_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3911_ _2121_/X _2201_/X _1994_/X _4336_/Q vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__o31a_1
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _3842_/A vssd1 vssd1 vccd1 vccd1 _4307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2722__B _4131_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3773_ _4272_/Q _3767_/X _3771_/X input87/X _3772_/X vssd1 vssd1 vccd1 vccd1 _4272_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2936__A1 _4041_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ _2726_/A _4132_/Q vssd1 vssd1 vccd1 vccd1 _2725_/A sky130_fd_sc_hd__and2_1
X_2655_ _3882_/C _4044_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _3271_/B sky130_fd_sc_hd__mux2_4
XANTENNA__3834__A _3847_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2586_ _2481_/X _2501_/X _2429_/X _2430_/X _4381_/Q vssd1 vssd1 vccd1 vccd1 _2586_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4325_ _4346_/CLK _4325_/D vssd1 vssd1 vccd1 vccd1 _4325_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2164__A2 _2160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__A3 _1998_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4284_/CLK _4256_/D vssd1 vssd1 vccd1 vccd1 _4256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4187_ _4225_/CLK _4187_/D vssd1 vssd1 vccd1 vccd1 _4187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4087__D _4087_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3207_ _3692_/A vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3138_ _3257_/B _4212_/Q _3144_/S vssd1 vssd1 vccd1 vccd1 _3646_/C sky130_fd_sc_hd__mux2_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3069_ _3208_/C _4193_/Q _3076_/S vssd1 vssd1 vccd1 vccd1 _3600_/A sky130_fd_sc_hd__mux2_2
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2624__B1 _2623_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2913__A _2913_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2927__A1 _4109_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3447__C _4002_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4080__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3352__A1 _3942_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2155__A2 _1971_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2312__C1 _4360_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2863__A0 _3843_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2615__B1 _2298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2823__A _2828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3919__A _3919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__B _3661_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output296_A _2908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__C1 _4365_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2440_ _2507_/A _3677_/A _2507_/C _2440_/D vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3654__A _3654_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2052__B1_N _4074_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2371_ _3532_/B _2362_/X _2364_/Y _2370_/Y vssd1 vssd1 vccd1 vccd1 _3963_/A sky130_fd_sc_hd__o211ai_4
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4250_/CLK _4110_/D vssd1 vssd1 vccd1 vccd1 _4110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _4051_/CLK _4041_/D vssd1 vssd1 vccd1 vccd1 _4041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2436__C _2436_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2606__B1 _2517_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2733__A _2737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2082__A1 _4351_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3829__A _3847_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4370__D _4370_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2909__A1 input52/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3825_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3845_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3756_ _4262_/Q _3750_/X _3754_/X _2466_/D _3755_/X vssd1 vssd1 vccd1 vccd1 _4262_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3267__C _3276_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2707_ _2715_/A _4124_/Q vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__and2_1
X_3687_ _3687_/A vssd1 vssd1 vccd1 vccd1 _4229_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3564__A _3564_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput242 _3156_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[1] sky130_fd_sc_hd__buf_2
Xoutput220 _3045_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput253 _2719_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[15] sky130_fd_sc_hd__buf_2
Xoutput231 _3050_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[2] sky130_fd_sc_hd__buf_2
X_2638_ _2638_/A _2638_/B _2638_/C _2638_/D vssd1 vssd1 vccd1 vccd1 _2638_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3334__A1 _4068_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3283__B _3283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput275 _2695_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[6] sky130_fd_sc_hd__buf_2
Xoutput264 _2741_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput286 _2853_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__3714__D _3724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2569_ _2281_/X _2566_/Y _2293_/X _2567_/Y _2568_/Y vssd1 vssd1 vccd1 vccd1 _2569_/Y
+ sky130_fd_sc_hd__o221ai_4
Xoutput297 _2913_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_88_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2542__C1 _2409_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4308_ _4371_/CLK _4308_/D vssd1 vssd1 vccd1 vccd1 _4308_/Q sky130_fd_sc_hd__dfxtp_1
X_4239_ _4264_/CLK _4239_/D vssd1 vssd1 vccd1 vccd1 _4239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4395__A _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3098__A0 _3227_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2908__A _2908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2845__A0 _3837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2643__A _3428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2073__A1 _4348_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4280__D _4280_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2081__C _2081_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2789__S _2825_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3474__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3325__A1 _4065_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input55_A cpu_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2818__A _2828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output211_A _3082_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output309_A _2807_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3649__A _3649_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ _4357_/Q vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__2064__A1 _4075_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2272__B _2272_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4190__D _4190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3610_ _3610_/A vssd1 vssd1 vccd1 vccd1 _4197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3541_ _3546_/A _3541_/B vssd1 vssd1 vccd1 vccd1 _4159_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3995__B1_N _2602_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3384__A _3384_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3472_ _2739_/A _2248_/X _3298_/A vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__2119__A2 _2257_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3815__C _3815_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3316__A1 _4059_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2423_ _2423_/A vssd1 vssd1 vccd1 vccd1 _2919_/A sky130_fd_sc_hd__buf_2
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2354_ _2514_/A vssd1 vssd1 vccd1 vccd1 _2644_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3831__B _3845_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2728__A _2739_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2285_ _2531_/A vssd1 vssd1 vccd1 vccd1 _2286_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4319__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2827__A0 _3215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4024_ _4085_/CLK _4024_/D vssd1 vssd1 vccd1 vccd1 _4024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4365__D _4365_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2182__B _2182_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3808_ _3808_/A vssd1 vssd1 vccd1 vccd1 _4293_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3555__B2 _2583_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3555__A1 _4170_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2358__A2 _2357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3739_ _4252_/Q _3734_/X _3735_/X input85/X _3738_/X vssd1 vssd1 vccd1 vccd1 _4252_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3294__A _3315_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2638__A _2638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2357__B _2357_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4275__D _4275_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3491__B1 _3489_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2076__C _2158_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3469__A _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2373__A _2469_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2046__A1 _2204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2597__A2 _2596_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2092__B _2207_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3188__B _3199_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3916__B _3916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3635__C _3635_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__D1 _2380_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output161_A _2603_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output259_A _2730_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2521__A2 _2366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__C _3370_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2070_ _3346_/A _3346_/B _2060_/Y _2064_/Y _2069_/Y vssd1 vssd1 vccd1 vccd1 _2085_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__2809__A0 _3821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4185__D _4185_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3379__A _3379_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_11_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2972_ _3036_/A vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2283__A _3441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2588__A2 _2582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _1923_/A vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_26_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3826__B _3845_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3524_ _3544_/A vssd1 vssd1 vccd1 vccd1 _3524_/X sky130_fd_sc_hd__buf_2
XANTENNA__4003__A _4003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3455_ _3455_/A _3459_/B _3455_/C vssd1 vssd1 vccd1 vccd1 _3456_/A sky130_fd_sc_hd__and3_1
XANTENNA__4141__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2406_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3842__A _3842_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3386_ _3386_/A _3405_/B _3400_/C vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__and3_1
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _2412_/A _2520_/B _2520_/C _2337_/D vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__nand4_2
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2268_ _4251_/Q vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2608__D _2608_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2276__A1 _2268_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4095__D _4095_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2892__S _2905_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4007_ _4085_/CLK _4007_/D vssd1 vssd1 vccd1 vccd1 _4007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4291__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2199_ _3343_/C vssd1 vssd1 vccd1 vccd1 _2200_/A sky130_fd_sc_hd__buf_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3289__A _3289_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2193__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3776__B2 input89/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3776__A1 _4274_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3455__C _3455_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3174__D _3190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3752__A _3769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2368__A _2575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3190__C _3195_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A cpu_adr_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3199__A _3221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2019__A1 _1993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4014__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3519__A1 _3730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3646__B _3659_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3138__S _3144_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3365__C _3365_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__D1 _3331_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3662__A _3662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3240_ _3240_/A vssd1 vssd1 vccd1 vccd1 _4031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3381__B _3381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3171_ _3591_/A vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _1942_/B _1971_/D _1971_/C _2121_/X vssd1 vssd1 vccd1 vccd1 _3945_/C sky130_fd_sc_hd__a31o_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2053_ _2053_/A _2074_/D _2053_/C _2072_/B vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__nand4_4
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3758__A1 _3752_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2955_ _3178_/C _4079_/Q _2955_/S vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3837__A _3837_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2741__A _2741_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2886_ _3853_/C _4032_/Q _2886_/S vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__mux2_4
XANTENNA__3556__B _3556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3048__S _3076_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2194__B1 _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3507_ _3510_/A _4139_/Q _3657_/C vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__and3_1
XANTENNA__2887__S _2911_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3930__A1 _2155_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3572__A _3586_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3438_ _3438_/A vssd1 vssd1 vccd1 vccd1 _4110_/D sky130_fd_sc_hd__clkbuf_1
X_3369_ _3369_/A vssd1 vssd1 vccd1 vccd1 _3389_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2497__A1 _2427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2188__A _2188_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3291__B _3689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2497__B2 _2430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4037__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3749__A1 _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3747__A _3764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4187__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2651__A _2896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3466__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3906__D1 _3938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2185__B1 _2184_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__A1 _4341_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3482__A _3876_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2797__S _2845_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput120 spi_dat_i[1] vssd1 vssd1 vccd1 vccd1 _3526_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2488__A1 _2486_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2098__A _2098_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput131 spi_dat_i[2] vssd1 vssd1 vccd1 vccd1 _2310_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput142 spi_rty_i vssd1 vssd1 vccd1 vccd1 _2383_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3988__A1 _3952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1999__B1 _1998_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3657__A _3657_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2740_ _2748_/A _4139_/Q vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__and2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2963__A2 _2200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2671_ _3276_/B _4116_/Q _2942_/S vssd1 vssd1 vccd1 vccd1 _3453_/C sky130_fd_sc_hd__mux2_4
XANTENNA__3376__B _3381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3343__D_N _2069_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2176__B1 _4347_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3392__A _3392_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3912__A1 _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4341_ _4346_/CLK _4341_/D vssd1 vssd1 vccd1 vccd1 _4341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4272_ _4280_/CLK _4272_/D vssd1 vssd1 vccd1 vccd1 _4272_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3823__C _3823_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2479__A1 _3541_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3223_ _3343_/B vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ _2972_/X _2974_/X _3569_/A vssd1 vssd1 vccd1 vccd1 _3154_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2158__D _2158_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2736__A _2736_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2105_ _4391_/Q vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__clkinv_2
X_3085_ _3217_/C _4197_/Q _3112_/S vssd1 vssd1 vccd1 vccd1 _3609_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3979__A1 _4371_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2036_ _4067_/Q vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2100__B1 _2099_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4373__D _4373_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _3968_/X _3969_/X _2559_/X _2563_/Y vssd1 vssd1 vccd1 vccd1 _4378_/D sky130_fd_sc_hd__o22a_1
XFILLER_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ _2943_/A _3447_/B _3439_/A vssd1 vssd1 vccd1 vccd1 _2939_/A sky130_fd_sc_hd__and3_1
XANTENNA__2403__A1 _2380_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2403__B2 _2509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3286__B _3689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3717__D _3724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2869_ _3845_/A _4029_/Q _2905_/S vssd1 vssd1 vccd1 vccd1 _3234_/C sky130_fd_sc_hd__mux2_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__D _4283_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2642__A1 _2328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3477__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2381__A _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input85_A gpio_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2812__C _3386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4202__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output241_A _3154_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3940__A _3940_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2556__A _4271_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2881__A1 _4031_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4352__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2275__B _2590_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4193__D _4193_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2633__A1 _2328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3910_ _4335_/Q _3908_/X _1983_/Y _3909_/X _3903_/X vssd1 vssd1 vccd1 vccd1 _4335_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _3841_/A _3845_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__and3_1
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3387__A _3387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2723_ _2723_/A vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2397__B1 _2396_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2654_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2950_/S sky130_fd_sc_hd__buf_2
XANTENNA__2149__B1 _2083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2585_ _4274_/Q _2295_/X _2298_/X input89/X vssd1 vssd1 vccd1 vccd1 _2585_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__3834__B _3853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4324_ _4326_/CLK _4324_/D vssd1 vssd1 vccd1 vccd1 _4324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4368__D _4368_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4255_ _4286_/CLK _4255_/D vssd1 vssd1 vccd1 vccd1 _4255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3850__A _3850_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3206_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3692_/A sky130_fd_sc_hd__clkbuf_4
X_4186_ _4284_/CLK _4186_/D vssd1 vssd1 vccd1 vccd1 _4186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3137_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3151_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2321__B1 _2320_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2466__A _2507_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3068_ _3068_/A vssd1 vssd1 vccd1 vccd1 _3068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2624__A1 _2622_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _1993_/X _2018_/X _4063_/Q vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__o21ai_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3297__A _3297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4225__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3352__A2 _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2155__A3 _1998_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4278__D _4278_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4375__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2376__A _2406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2312__B1 _2311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2863__A1 _4028_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2615__A1 _4278_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2615__B2 input93/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2823__B _2841_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__C _3648_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_2_1_0_CLK_A clkbuf_2_1_0_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3000__A _3000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__B1 _2377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output191_A _3020_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output289_A _2873_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__A _3935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4188__D _4188_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2551__B1 _2298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2370_ _2262_/X _2375_/A _2408_/A _2409_/A _2369_/Y vssd1 vssd1 vccd1 vccd1 _2370_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__3670__A _3670_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ _4380_/CLK _4040_/D vssd1 vssd1 vccd1 vccd1 _4040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2286__A _2286_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2436__D _2503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2606__B2 _2450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2606__A1 _2427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3829__B _3829_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2733__B _4136_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2082__A2 _2182_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4248__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3824_ _3824_/A vssd1 vssd1 vccd1 vccd1 _4300_/D sky130_fd_sc_hd__clkbuf_1
X_3755_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3567__C1 _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3267__D _3271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2706_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__clkbuf_1
X_3686_ _3699_/A _4229_/Q _3703_/C _3689_/D vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__and4_1
XANTENNA__3845__A _3845_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput210 _3078_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[10] sky130_fd_sc_hd__buf_2
X_2637_ _4281_/Q vssd1 vssd1 vccd1 vccd1 _2637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3564__B _3564_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2790__A0 _3815_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3319__C1 _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput221 _3114_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput232 _3149_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput243 _3158_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__3056__S _3076_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3334__A2 _3331_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3283__C _3323_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput265 _2743_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput254 _2721_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput276 _2699_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[7] sky130_fd_sc_hd__buf_2
X_2568_ _2301_/X _2302_/X _2324_/X _2552_/X _4379_/Q vssd1 vssd1 vccd1 vccd1 _2568_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2542__B1 _2408_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput298 _2918_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput287 _2860_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__4098__D _4098_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2499_ _2499_/A vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3580__A _3580_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _4371_/CLK _4307_/D vssd1 vssd1 vccd1 vccd1 _4307_/Q sky130_fd_sc_hd__dfxtp_1
X_4238_ _4264_/CLK _4238_/D vssd1 vssd1 vccd1 vccd1 _4238_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3098__A1 _4201_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2196__A _3023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4169_ _4180_/CLK _4169_/D vssd1 vssd1 vccd1 vccd1 _4169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2845__A1 _4025_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2924__A _2924_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2073__A2 _2012_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2135__S _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3755__A _3772_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2081__D _2081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3474__B _4123_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3325__A2 _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input48_A cpu_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3490__A _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2818__B _2841_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output204_A _2982_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2834__A _2859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2064__A2 _2152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _2462_/C _3536_/X _3528_/X _2463_/Y _3537_/X vssd1 vssd1 vccd1 vccd1 _4158_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3665__A _3665_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2772__A0 _3188_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3471_ _4122_/Q _3350_/X _4395_/A _3469_/X _3470_/X vssd1 vssd1 vccd1 vccd1 _4122_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2422_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2423_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3316__A2 _3314_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2353_ _4152_/Q vssd1 vssd1 vccd1 vccd1 _2353_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3831__C _3831_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2284_ _2284_/A vssd1 vssd1 vccd1 vccd1 _2531_/A sky130_fd_sc_hd__buf_4
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4023_ _4051_/CLK _4023_/D vssd1 vssd1 vccd1 vccd1 _4023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2827__A1 _4092_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2744__A _2748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3788__C1 _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4070__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4381__D _4381_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2460__C1 _2373_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ _3807_/A _3821_/B _3903_/A vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__and3_1
XANTENNA__3555__A2 _3447_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3575__A _3575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1999_ _4332_/Q _2182_/B _1998_/Y _1973_/X _1965_/X vssd1 vssd1 vccd1 vccd1 _3294_/B
+ sky130_fd_sc_hd__o2111ai_4
X_3738_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3294__B _3294_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2763__A0 _4292_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3669_ _3798_/A _3673_/B _3669_/C vssd1 vssd1 vccd1 vccd1 _3670_/A sky130_fd_sc_hd__or3_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2919__A _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__B _2638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2357__C _2357_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2279__C1 _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3491__A1 _4130_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3491__B2 _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2654__A _2898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input102_A gpio_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3779__C1 _3774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2046__A2 _2018_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4291__D _4291_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2451__C1 _4368_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3188__C _3188_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3485__A _3976_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3916__C _3916_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__C1 _3800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2829__A _2829_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output154_A _2555_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2634__B1_N _4177_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2809__A1 _4019_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4093__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _2197_/X _2200_/X _3667_/A vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__o21a_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _4356_/Q vssd1 vssd1 vccd1 vccd1 _2201_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3395__A _3395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3826__C _3831_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3523_ _3536_/A vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__clkbuf_4
X_3454_ _3454_/A vssd1 vssd1 vccd1 vccd1 _4116_/D sky130_fd_sc_hd__clkbuf_1
X_2405_ _2379_/X _2399_/Y _2404_/X _2373_/X vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__o211a_2
XANTENNA__2739__A _2739_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3385_ _3433_/A vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2336_ _2336_/A vssd1 vssd1 vccd1 vccd1 _2520_/C sky130_fd_sc_hd__buf_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2267_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2409_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4376__D _4376_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4006_ _4391_/Q _2357_/A _3953_/B _3953_/A _3938_/D vssd1 vssd1 vccd1 vccd1 _4391_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__2474__A _2474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2276__A2 _2539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2198_ _2349_/A vssd1 vssd1 vccd1 vccd1 _3343_/C sky130_fd_sc_hd__buf_2
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3776__A2 _3767_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2433__C1 _2373_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2984__B1 _3675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3933__C1 _3912_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2368__B _2520_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4286__D _4286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3190__D _3190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2384__A _2384_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3199__B _3199_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2019__A2 _2018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2975__A0 _3283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3646__C _3646_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3519__A2 _2428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4309__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output271_A _2753_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__C1 _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3943__A _3943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3381__C _3400_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3170_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__buf_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4196__D _4196_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2121_ _2121_/A vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__buf_2
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2052_ _2136_/A _2015_/X _4074_/Q vssd1 vssd1 vccd1 vccd1 _3346_/A sky130_fd_sc_hd__a21boi_1
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2294__A _3578_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3758__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2966__A0 _3273_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3837__B _3845_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2954_ _3796_/A _4009_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _3178_/C sky130_fd_sc_hd__mux2_2
X_2885_ _4312_/Q input48/X _2885_/S vssd1 vssd1 vccd1 vccd1 _3853_/C sky130_fd_sc_hd__mux2_2
XANTENNA__2194__A1 _2128_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3506_ _3976_/A vssd1 vssd1 vccd1 vccd1 _3657_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3853__A _3871_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3572__B _3586_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3930__A2 _2072_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3437_ _3457_/A _3437_/B _3437_/C vssd1 vssd1 vccd1 vccd1 _3438_/A sky130_fd_sc_hd__or3_1
XANTENNA__2469__A _2469_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2497__A2 _2428_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3368_ _3368_/A vssd1 vssd1 vccd1 vccd1 _4081_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3291__C _3291_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2188__B _2211_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2319_ _2529_/A vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__buf_2
XFILLER_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3343_/A _3326_/C _3323_/C _1990_/Y vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__or4b_1
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3749__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2957__A0 _4290_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3466__C _3466_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3906__C1 _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2185__A1 _4065_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__A2 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__A0 _3253_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput110 spi_dat_i[10] vssd1 vssd1 vccd1 vccd1 _2448_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2488__A2 _2411_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2098__B _2098_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput132 spi_dat_i[30] vssd1 vssd1 vccd1 vccd1 _2635_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput121 spi_dat_i[20] vssd1 vssd1 vccd1 vccd1 _2561_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input30_A cpu_adr_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3988__A2 _3955_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3003__A _3003_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1999__A1 _4332_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2842__A _2842_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3938__A _3938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2948__B1 _3354_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4131__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _3657_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3376__C _3376_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2670_ _3887_/C _4046_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__mux2_4
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4281__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3673__A _3798_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2176__A1 _2121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3912__A2 _1996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4340_ _4347_/CLK _4340_/D vssd1 vssd1 vccd1 vccd1 _4340_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2289__A _2387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4271_ _4275_/CLK _4271_/D vssd1 vssd1 vccd1 vccd1 _4271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _3222_/A vssd1 vssd1 vccd1 vccd1 _4025_/D sky130_fd_sc_hd__clkbuf_1
X_3153_ _3167_/C _4181_/Q _3157_/S vssd1 vssd1 vccd1 vccd1 _3569_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2479__A2 _2362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2104_ _3696_/A vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__buf_2
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1921__A _1938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3084_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3112_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__C1 _4388_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3979__A2 _3965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2035_ _2032_/Y _1962_/A _2034_/Y vssd1 vssd1 vccd1 vccd1 _3326_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__2100__A1 _2106_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3848__A _3848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2752__A _2752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3986_ _3952_/X _3955_/X _2554_/Y vssd1 vssd1 vccd1 vccd1 _4377_/D sky130_fd_sc_hd__o21bai_1
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2403__A2 _3564_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2937_ _3265_/C _4111_/Q _2937_/S vssd1 vssd1 vccd1 vccd1 _3439_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3059__S _3073_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3286__C _3286_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2868_ _4309_/Q input44/X _2904_/S vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__mux2_8
X_2799_ _2799_/A _2812_/B _3381_/A vssd1 vssd1 vccd1 vccd1 _2800_/A sky130_fd_sc_hd__and3_2
XANTENNA__3583__A _3583_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3116__A0 _3241_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2199__A _3343_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4154__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2627__C1 _2246_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__A2 _2329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2662__A _2662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3477__B _4125_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3493__A _3493_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input78_A gpio_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3940__B _3942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output234_A _3053_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2618__C1 _2579_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2275__C _2414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2633__A2 _2329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3668__A _3668_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2094__B1 _1986_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _3840_/A vssd1 vssd1 vccd1 vccd1 _4306_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3310__D_N _2207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3771_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2722_ _2726_/A _4131_/Q vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__and2_1
XANTENNA__2397__A1 _2390_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2653_ _2662_/A vssd1 vssd1 vccd1 vccd1 _2898_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2149__A1 _2662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2584_ _3466_/C _4170_/Q _2583_/X _3544_/A vssd1 vssd1 vccd1 vccd1 _2584_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__3834__C _3834_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4027__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4323_ _4356_/CLK _4323_/D vssd1 vssd1 vccd1 vccd1 _4323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4284_/CLK _4254_/D vssd1 vssd1 vccd1 vccd1 _4254_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3850__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2747__A _2747_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4177__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2321__A1 _3529_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4185_ _4225_/CLK _4185_/D vssd1 vssd1 vccd1 vccd1 _4185_/Q sky130_fd_sc_hd__dfxtp_1
X_3205_ _3205_/A vssd1 vssd1 vccd1 vccd1 _4018_/D sky130_fd_sc_hd__clkbuf_1
X_3136_ _3136_/A vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2466__B _3677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3067_ _3081_/A _3070_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _3068_/A sky130_fd_sc_hd__and3_1
XANTENNA__4384__D _4384_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2071__A1_N _4068_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2018_ _2018_/A vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3578__A _3578_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2624__A2 _2366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2388__A1 _2386_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3969_ _3992_/A vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2560__A1 _2386_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input132_A spi_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2312__A1 _2256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2312__B2 _2260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4294__D _4294_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3488__A _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2615__A2 _2322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2392__A _2412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2823__C _3391_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2379__A1 _2375_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__B2 _3769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output184_A _3007_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__B _3935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2000__B1 _4053_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2551__A1 _4270_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2551__B2 input84/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2606__A2 _2449_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2067__B1 _2066_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3398__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3829__C _3829_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3823_ _3823_/A _3829_/B _3823_/C vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__or3_1
XANTENNA__3567__B1 _2407_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3754_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2705_ _2705_/A vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__clkbuf_1
X_3685_ _3707_/A vssd1 vssd1 vccd1 vccd1 _3703_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3845__B _3845_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput200 _3037_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[31] sky130_fd_sc_hd__buf_2
X_2636_ _2427_/A _2428_/A _2517_/X _2434_/A _4388_/Q vssd1 vssd1 vccd1 vccd1 _2636_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2790__A1 _4016_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3319__B1 _2165_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput211 _3082_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput233 _3152_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput222 _3118_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput244 _3160_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__4379__D _4379_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput255 _2723_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[17] sky130_fd_sc_hd__buf_2
Xoutput277 _2703_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput266 _2745_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[27] sky130_fd_sc_hd__buf_2
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2567_ _4272_/Q _2322_/X _2298_/A input87/X vssd1 vssd1 vccd1 vccd1 _2567_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__2542__A1 _2406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3861__A _3861_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3283__D _3317_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput299 _2924_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput288 _2867_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2498_ _2419_/X _3543_/B _2497_/Y vssd1 vssd1 vccd1 vccd1 _2498_/Y sky130_fd_sc_hd__o21ai_1
X_4306_ _4371_/CLK _4306_/D vssd1 vssd1 vccd1 vccd1 _4306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4237_ _4264_/CLK _4237_/D vssd1 vssd1 vccd1 vccd1 _4237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3580__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4168_ _4172_/CLK _4168_/D vssd1 vssd1 vccd1 vccd1 _4168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3119_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4099_ _4286_/CLK _4099_/D vssd1 vssd1 vccd1 vccd1 _4099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2058__B1 _4353_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3101__A _3137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2230__B1 _2138_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3474__C _4002_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4342__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4289__D _4289_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3771__A _3771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2387__A _2387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2818__C _3389_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3494__C1 _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2834__B _2841_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3011__A _3011_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3946__A _3946_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3157__S _3157_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2772__A1 _4083_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3470_ _3470_/A vssd1 vssd1 vccd1 vccd1 _3470_/X sky130_fd_sc_hd__buf_2
XANTENNA__4199__D _4199_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3681__A _3699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2421_ _2421_/A vssd1 vssd1 vccd1 vccd1 _2421_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2352_ _2700_/A _2678_/A _2248_/X _2286_/A _2352_/D1 vssd1 vssd1 vccd1 vccd1 _2356_/A
+ sky130_fd_sc_hd__o2111ai_4
X_2283_ _3441_/A vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2297__A _2533_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4022_ _4085_/CLK _4022_/D vssd1 vssd1 vccd1 vccd1 _4022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2744__B _4141_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4215__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3788__B1 _2407_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2460__B1 _3973_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3856__A _3856_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4365__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _4292_/D sky130_fd_sc_hd__clkbuf_1
X_3737_ _3765_/A _3736_/Y _3264_/A vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__o21ai_4
X_1998_ input32/X _1998_/B _2053_/A _2081_/D vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3294__C _3294_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2763__A1 input46/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3668_ _3668_/A vssd1 vssd1 vccd1 vccd1 _4221_/D sky130_fd_sc_hd__clkbuf_1
X_2619_ _2423_/A _2387_/A _4175_/Q vssd1 vssd1 vccd1 vccd1 _2619_/Y sky130_fd_sc_hd__a21boi_1
X_3599_ _3599_/A vssd1 vssd1 vccd1 vccd1 _4192_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3591__A _3591_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2515__A1 _2330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2638__C _2638_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3476__C1 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2279__B1 _2246_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3491__A2 _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3779__B1 _2609_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2451__B1 _2311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3188__D _3208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2203__B1 _2202_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3916__D _3938_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__B1 _3945_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input60_A cpu_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3006__A _3010_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output147_A _2480_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4238__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output314_A _2956_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2690__A0 _3286_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2970_ _3279_/C _4221_/Q _3335_/A vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2442__B1 _2441_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ _1938_/A vssd1 vssd1 vccd1 vccd1 _2184_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3676__A _3676_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3522_ _3564_/B _3522_/B vssd1 vssd1 vccd1 vccd1 _4147_/D sky130_fd_sc_hd__nor2_1
X_3453_ _3457_/A _3462_/B _3453_/C vssd1 vssd1 vccd1 vccd1 _3454_/A sky130_fd_sc_hd__or3_1
X_2404_ _2499_/A vssd1 vssd1 vccd1 vccd1 _2404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1924__A _1924_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3384_ _3384_/A vssd1 vssd1 vccd1 vccd1 _4088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2335_ _2335_/A vssd1 vssd1 vccd1 vccd1 _2520_/B sky130_fd_sc_hd__buf_2
X_2266_ _2367_/A _2335_/A _2117_/X vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__a21o_2
X_2197_ _3036_/A vssd1 vssd1 vccd1 vccd1 _2197_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ _3991_/A _3992_/A _2224_/X _2245_/X vssd1 vssd1 vccd1 vccd1 _4390_/D sky130_fd_sc_hd__o22a_1
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2755__A _2957_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__A0 _4328_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2433__B1 _2404_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2984__A1 _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3586__A _3586_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3933__B1 _3932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2368__C _2520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2665__A _2683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2672__B1 _3453_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3199__C _3199_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3496__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2975__A1 _4222_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4346_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3924__B1 _2179_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output264_A _2741_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3688__C1 _3683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4060__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2120_ _2120_/A vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2575__A _2575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2051_ _3326_/B _3328_/A _2051_/C vssd1 vssd1 vccd1 vccd1 _2085_/B sky130_fd_sc_hd__nor3_1
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3758__A3 _3748_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2953_ _4289_/Q input69/X _2953_/S vssd1 vssd1 vccd1 vccd1 _3796_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2966__A1 _4219_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ _2884_/A vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3837__C _3855_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2194__A2 _2133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3505_ _4138_/Q _3488_/X _3489_/X _3490_/X _3504_/X vssd1 vssd1 vccd1 vccd1 _4138_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3853__B _3853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3572__C _3572_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__C1 _3504_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3436_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4387__D _4387_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3367_ _3367_/A _3381_/B _3376_/C vssd1 vssd1 vccd1 vccd1 _3368_/A sky130_fd_sc_hd__and3_1
XANTENNA__3291__D _3925_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2188__C _2211_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2351__C1 _2350_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2318_ _2224_/X _2245_/X _3957_/A _2125_/X vssd1 vssd1 vccd1 vccd1 _2318_/X sky130_fd_sc_hd__o211a_2
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3298_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3326_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2249_ _2382_/A _2383_/A _2384_/A vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__nor3b_1
XANTENNA__3080__S _3109_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3749__A3 _3748_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2957__A1 input70/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3906__B1 _1988_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4083__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2185__A2 _1977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__A1 _4211_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput100 gpio_dat_i[4] vssd1 vssd1 vccd1 vccd1 _2337_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput111 spi_dat_i[11] vssd1 vssd1 vccd1 vccd1 _2462_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4297__D _4297_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput133 spi_dat_i[31] vssd1 vssd1 vccd1 vccd1 _2644_/C sky130_fd_sc_hd__clkbuf_2
Xinput122 spi_dat_i[21] vssd1 vssd1 vccd1 vccd1 _3553_/A1 sky130_fd_sc_hd__buf_2
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2893__A0 _3243_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2098__C _2098_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input23_A cpu_adr_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2395__A _2414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2645__B1 _2644_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1999__A2 _2182_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3938__B _3938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2948__A1 _2677_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3657__C _3657_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3954__A _3954_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3673__B _3673_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2176__A2 _2160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4270_ _4282_/CLK _4270_/D vssd1 vssd1 vccd1 vccd1 _4270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3221_ _3221_/A _3227_/B _3221_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _3222_/A sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_9_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4141_/CLK sky130_fd_sc_hd__clkbuf_16
X_3152_ _3152_/A vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2333__C1 _4362_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2103_ _2590_/A vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3083_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2636__B1 _2517_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2034_ input16/X _2168_/A _2033_/Y _1938_/A vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2100__A2 _2112_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2752__B _4145_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3985_ _3968_/X _3969_/X _2542_/X _2547_/Y vssd1 vssd1 vccd1 vccd1 _4376_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _3874_/A _4041_/Q _2936_/S vssd1 vssd1 vccd1 vccd1 _3265_/C sky130_fd_sc_hd__mux2_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2867_ _2867_/A vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3286__D _3286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3864__A _3864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3993__B1_N _2587_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2798_ _3199_/C _4087_/Q _2955_/S vssd1 vssd1 vccd1 vccd1 _3381_/A sky130_fd_sc_hd__mux2_2
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3419_ _3419_/A vssd1 vssd1 vccd1 vccd1 _4102_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3116__A1 _4206_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2875__A0 _4310_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3104__A _3104_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2627__B1 _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2943__A _2943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3477__C _4002_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3774__A _3774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3940__C _3940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output227_A _3136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3014__A _3014_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2618__B1 _2617_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2079__D1 _1985_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2853__A _2853_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2275__D _2275_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3949__A _3949_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2094__A1 _1976_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3043__A0 _3186_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3770_ _3769_/X _3764_/X _3765_/X _2558_/Y _3757_/X vssd1 vssd1 vccd1 vccd1 _4271_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2721_ _2721_/A vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2397__A2 _3673_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2149__A2 _2148_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ _4324_/Q input2/X _2949_/S vssd1 vssd1 vccd1 vccd1 _3882_/C sky130_fd_sc_hd__mux2_2
X_2583_ _2628_/A _2644_/B _2583_/C vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__and3_1
XFILLER_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2554__C1 _2553_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4322_ _4391_/CLK _4322_/D vssd1 vssd1 vccd1 vccd1 _4322_/Q sky130_fd_sc_hd__dfxtp_1
X_4253_ _4284_/CLK _4253_/D vssd1 vssd1 vccd1 vccd1 _4253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2306__C1 _2305_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3204_ _3224_/A _3204_/B _3224_/C _3219_/D vssd1 vssd1 vccd1 vccd1 _3205_/A sky130_fd_sc_hd__or4_1
XANTENNA__1932__A _2007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4184_ _4262_/CLK _4184_/D vssd1 vssd1 vccd1 vccd1 _4184_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3850__C _3855_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2857__A0 _3841_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3135_ _3135_/A _3142_/B _3644_/A vssd1 vssd1 vccd1 vccd1 _3136_/A sky130_fd_sc_hd__and3_1
XANTENNA__2321__A2 _2283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2466__C _2507_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2609__B1 _2608_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3066_ _3204_/B _4192_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3598_/C sky130_fd_sc_hd__mux2_1
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3859__A _3859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2017_ _1962_/A _2012_/Y _2013_/Y _2016_/Y vssd1 vssd1 vccd1 vccd1 _3320_/B sky130_fd_sc_hd__a31oi_4
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3968_ _3991_/A vssd1 vssd1 vccd1 vccd1 _3968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2388__A2 _3468_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2919_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3594__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3899_ _3899_/A vssd1 vssd1 vccd1 vccd1 _4331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2560__A2 _2424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2938__A _2943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2312__A2 _2258_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input125_A spi_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3769__A _3769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4271__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input90_A gpio_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__A2 _2376_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3935__C _3935_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3009__A _3009_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output177_A _2992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__C1 _2535_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2000__A1 _1993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2551__A2 _2322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2848__A _2848_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2839__A0 _3834_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2583__A _2628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2067__A1 _2065_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3398__B _3413_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3822_ _3822_/A vssd1 vssd1 vccd1 vccd1 _4299_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3567__A1 _4180_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3753_ _3752_/X _3747_/X _3748_/X _2457_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _4261_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__1927__A _2011_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2704_ _2704_/A _4123_/Q vssd1 vssd1 vccd1 vccd1 _2705_/A sky130_fd_sc_hd__and2_1
X_3684_ _4228_/Q _3351_/X _4394_/A _3678_/X _3683_/X vssd1 vssd1 vccd1 vccd1 _4228_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3845__C _3855_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput201 _2971_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[3] sky130_fd_sc_hd__buf_2
X_2635_ _2635_/A1 _2628_/A _2514_/X _2531_/A _2634_/Y vssd1 vssd1 vccd1 vccd1 _3562_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__3319__A1 _4061_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput223 _3123_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput212 _3087_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput234 _3053_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__4144__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput267 _2747_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[28] sky130_fd_sc_hd__buf_2
Xoutput256 _2725_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput245 _4394_/X vssd1 vssd1 vccd1 vccd1 gpio_stb_o sky130_fd_sc_hd__buf_2
X_2566_ _3553_/A1 _2420_/X _2421_/X _2565_/Y vssd1 vssd1 vccd1 vccd1 _2566_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_88_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2542__A2 _2407_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3861__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4305_ _4356_/CLK _4305_/D vssd1 vssd1 vccd1 vccd1 _4305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput289 _2873_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput278 _2705_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2497_ _2427_/X _2428_/X _2303_/X _2430_/X _4372_/Q vssd1 vssd1 vccd1 vccd1 _2497_/Y
+ sky130_fd_sc_hd__o221ai_1
X_4236_ _4264_/CLK _4236_/D vssd1 vssd1 vccd1 vccd1 _4236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3580__C _3600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4294__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4177_/CLK _4167_/D vssd1 vssd1 vccd1 vccd1 _4167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3118_ _3118_/A vssd1 vssd1 vccd1 vccd1 _3118_/X sky130_fd_sc_hd__clkbuf_1
X_4098_ _4180_/CLK _4098_/D vssd1 vssd1 vccd1 vccd1 _4098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3589__A _3589_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3049_ _3063_/A _3052_/B _3584_/A vssd1 vssd1 vccd1 vccd1 _3050_/A sky130_fd_sc_hd__and3_1
XANTENNA__2058__A1 _1952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2230__A1 _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2518__C1 _4374_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3494__B1 _3489_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3499__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2834__C _3396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4017__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output294_A _2895_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4167__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2420_ _3441_/A vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__buf_2
XANTENNA__3681__B _4227_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2351_ _2343_/Y _3641_/A _2407_/A _2406_/A _2350_/Y vssd1 vssd1 vccd1 vccd1 _2357_/B
+ sky130_fd_sc_hd__o221ai_4
X_2282_ _2543_/A vssd1 vssd1 vccd1 vccd1 _3441_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4021_ _4051_/CLK _4021_/D vssd1 vssd1 vccd1 vccd1 _4021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3788__A1 _4285_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3788__B2 _2406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3202__A _3297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2460__A1 _2328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _1993_/X _1996_/X _4052_/Q vssd1 vssd1 vccd1 vccd1 _3294_/C sky130_fd_sc_hd__o21ai_1
X_3805_ _3823_/A _3805_/B _3805_/C vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__or3_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3736_ _2117_/X _2539_/A _2453_/A vssd1 vssd1 vccd1 vccd1 _3736_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3667_ _3667_/A _3796_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__and3_1
XANTENNA__3872__A _3872_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2618_ _2581_/X _2582_/X _2617_/Y _2579_/X vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__o211a_1
X_3598_ _3611_/A _3611_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__or3_1
XANTENNA__3323__D_N _2186_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2549_ _2319_/X _2289_/X _4166_/Q vssd1 vssd1 vccd1 vccd1 _2549_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__2515__A2 _2446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__D _2638_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4219_ _4225_/CLK _4219_/D vssd1 vssd1 vccd1 vccd1 _4219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3476__B1 _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2279__A1 _2224_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3779__A1 _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2309__B1_N _4149_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2451__B2 _2450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2451__A1 _2363_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2203__A1 _2201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3951__A1 _3728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input53_A cpu_dat_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2398__A _2509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3006__B _4235_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2690__A1 _4119_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3022__A _3022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output307_A _2793_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3957__A _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2861__A _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2442__B2 _2398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2442__A1 _2380_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ _1934_/A vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__buf_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ _3549_/A vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__buf_2
XANTENNA__3692__A _3692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3452_ _3452_/A vssd1 vssd1 vccd1 vccd1 _4115_/D sky130_fd_sc_hd__clkbuf_1
X_3383_ _3383_/A _3389_/B _3383_/C vssd1 vssd1 vccd1 vccd1 _3384_/A sky130_fd_sc_hd__or3_1
X_2403_ _2380_/A _3564_/A _2239_/Y _2509_/A _2402_/Y vssd1 vssd1 vccd1 vccd1 _2499_/A
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2101__A _2237_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2334_ _4255_/Q vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2408_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1940__A _4357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2196_ _3023_/A vssd1 vssd1 vccd1 vccd1 _3036_/A sky130_fd_sc_hd__buf_2
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4004_ _3991_/X _3992_/X _2648_/Y vssd1 vssd1 vccd1 vccd1 _4389_/D sky130_fd_sc_hd__o21bai_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4332__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__A1 input28/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3867__A _3871_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2433__A1 _2417_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2984__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3586__B _3586_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3719_ _4246_/Q _3167_/B _3044_/A _3697_/A _3705_/X vssd1 vssd1 vccd1 vccd1 _4246_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3933__A1 input20/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3107__A _3107_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2011__A _2011_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2368__D _2368_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2672__A1 _2128_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3199__D _3208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3496__B _4133_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3924__A1 _2044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4205__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3017__A _3021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3688__B1 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output257_A _2727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4355__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2856__A _2958_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2575__B _2638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2050_ _2050_/A _2050_/B _2050_/C _2050_/D vssd1 vssd1 vccd1 vccd1 _2051_/C sky130_fd_sc_hd__nand4_1
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _2704_/A _2133_/A _3358_/C vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3687__A _3687_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2883_ _2888_/A _2901_/B _3415_/A vssd1 vssd1 vccd1 vccd1 _2884_/A sky130_fd_sc_hd__and3_1
XANTENNA__2179__B1 _4344_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3504_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3504_/X sky130_fd_sc_hd__buf_2
XANTENNA__3853__C _3853_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1935__A _2059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3435_ _3435_/A vssd1 vssd1 vccd1 vccd1 _4109_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3679__B1 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3366_ _3366_/A vssd1 vssd1 vccd1 vccd1 _4080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2351__B1 _2407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2317_ _3527_/B _2255_/X _2312_/Y _2316_/Y vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__o211ai_4
X_3297_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3343_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2514_/A vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__buf_4
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2179_ _1952_/X _1932_/X _4344_/Q vssd1 vssd1 vccd1 vccd1 _2179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3597__A _3597_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2006__A input9/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4228__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3906__A1 _1987_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4378__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput101 gpio_dat_i[5] vssd1 vssd1 vccd1 vccd1 _3744_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput123 spi_dat_i[22] vssd1 vssd1 vccd1 vccd1 _2572_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput112 spi_dat_i[12] vssd1 vssd1 vccd1 vccd1 _2472_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput134 spi_dat_i[3] vssd1 vssd1 vccd1 vccd1 _3529_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2893__A1 _4103_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2098__D _2098_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2172__B1_N _4340_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A cpu_adr_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2645__B2 _2286_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2645__A1 _3444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3938__C _3938_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2948__A2 _2680_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3300__A _3300_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3673__C _3673_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3220_ _3220_/A vssd1 vssd1 vccd1 vccd1 _4024_/D sky130_fd_sc_hd__clkbuf_1
X_3151_ _3151_/A _3657_/B _3655_/C vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__and3_1
XANTENNA__2333__B1 _2311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _2638_/A vssd1 vssd1 vccd1 vccd1 _2590_/A sky130_fd_sc_hd__buf_2
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3082_ _3082_/A vssd1 vssd1 vccd1 vccd1 _3082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__A1 _2427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2636__B2 _2434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2097__C1 _2207_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2033_ _2120_/A _2141_/A _4346_/Q vssd1 vssd1 vccd1 vccd1 _2033_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _3952_/X _3955_/X _2536_/Y vssd1 vssd1 vccd1 vccd1 _4375_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__3210__A _3224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2935_ _4321_/Q input58/X _2935_/S vssd1 vssd1 vccd1 vccd1 _3874_/A sky130_fd_sc_hd__mux2_4
XFILLER_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2866_ _2888_/A _2872_/B _3407_/C vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__and3_1
X_2797_ _3817_/A _4017_/Q _2845_/S vssd1 vssd1 vccd1 vccd1 _3199_/C sky130_fd_sc_hd__mux2_2
XANTENNA__2572__B1 _2571_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3880__A _3880_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3418_ _3431_/A _3437_/B _3418_/C vssd1 vssd1 vccd1 vccd1 _3419_/A sky130_fd_sc_hd__or3_1
XFILLER_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3349_ _3724_/C vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input8_A cpu_adr_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2875__A1 input45/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2627__A1 _2581_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2943__B _3447_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3120__A _3120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4050__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2563__B1 _2562_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__C1 _3757_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3790__A _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4101__D _4101_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3512__C1 _3504_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2315__B1 _2314_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2618__A1 _2581_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2079__C1 _2137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3949__B _3973_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2094__A2 _2184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3030__A _3032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3043__A1 _4186_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _2726_/A _4130_/Q vssd1 vssd1 vccd1 vccd1 _2721_/A sky130_fd_sc_hd__and2_1
XANTENNA__3965__A _3965_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2651_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2949_/S sky130_fd_sc_hd__buf_2
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2554__B1 _2293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2582_ _2582_/A vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2003__C1 _1962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__C1 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4321_ _4371_/CLK _4321_/D vssd1 vssd1 vccd1 vccd1 _4321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4252_ _4284_/CLK _4252_/D vssd1 vssd1 vccd1 vccd1 _4252_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4011__D _4011_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2306__B1 _2293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3203_ _3343_/C vssd1 vssd1 vccd1 vccd1 _3224_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4183_ _4225_/CLK _4183_/D vssd1 vssd1 vccd1 vccd1 _4183_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3205__A _3205_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2857__A1 _4027_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2321__A3 _2286_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3134_ _3253_/C _4211_/Q _3147_/S vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2002__B1_N _4333_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3065_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3081_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2466__D _2466_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2609__A1 _2607_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4073__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2016_ _2136_/A _2015_/X _4062_/Q vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2490__C1 _2469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3967_ _4365_/Q _3965_/X _2399_/Y _3966_/Y vssd1 vssd1 vccd1 vccd1 _4365_/D sky130_fd_sc_hd__a211o_1
X_2918_ _2918_/A vssd1 vssd1 vccd1 vccd1 _2918_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2242__C1 _2264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3875__A _3875_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3594__B _3611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3898_ _3898_/A _3942_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__and3_1
X_2849_ _4306_/Q input41/X _2885_/S vssd1 vssd1 vccd1 vccd1 _3839_/C sky130_fd_sc_hd__mux2_2
XANTENNA__2545__B1 _2544_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3742__C1 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2938__B _3447_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3115__A _3115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input118_A spi_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3785__A _3945_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input83_A gpio_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2784__A0 _4295_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__C1 _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2536__B1 _2509_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3733__C1 _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2000__A2 _1996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3025__A _3025_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2839__A1 _4024_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4096__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2864__A _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2583__B _2644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2067__A2 _2001_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3398__C _3398_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3821_ _3821_/A _3821_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__and3_1
XANTENNA__3695__A _3695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3567__A2 _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2803__S _2826_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3752_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2703_ _2703_/A vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__clkbuf_1
X_3683_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2104__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2634_ _2423_/A _2387_/A _4177_/Q vssd1 vssd1 vccd1 vccd1 _2634_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__3319__A2 _3314_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput213 _3090_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput202 _2976_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput224 _3126_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput235 _3058_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[4] sky130_fd_sc_hd__buf_2
X_2565_ _2319_/X _2289_/X _4168_/Q vssd1 vssd1 vccd1 vccd1 _2565_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__2527__B1 _2387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput268 _2749_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[29] sky130_fd_sc_hd__buf_2
Xoutput257 _2727_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_99_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput246 _2217_/X vssd1 vssd1 vccd1 vccd1 gpio_we_o sky130_fd_sc_hd__buf_2
XANTENNA__3861__C _3879_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4304_ _4391_/CLK _4304_/D vssd1 vssd1 vccd1 vccd1 _4304_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1943__A _2001_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput279 _4395_/A vssd1 vssd1 vccd1 vccd1 spi_cyc_o sky130_fd_sc_hd__buf_2
X_2496_ _2496_/A1 _2420_/X _2421_/X _2495_/Y vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__a31oi_4
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4235_ _4264_/CLK _4235_/D vssd1 vssd1 vccd1 vccd1 _4235_/Q sky130_fd_sc_hd__dfxtp_1
X_4166_ _4172_/CLK _4166_/D vssd1 vssd1 vccd1 vccd1 _4166_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2571__B1_N _4169_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3117_/A _3125_/B _3631_/C vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__and3_1
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2774__A _2774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _4225_/CLK _4097_/D vssd1 vssd1 vccd1 vccd1 _4097_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3589__B _3609_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3048_ _3188_/C _4187_/Q _3076_/S vssd1 vssd1 vccd1 vccd1 _3584_/A sky130_fd_sc_hd__mux2_2
XANTENNA__2058__A2 _2160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2766__A0 _3186_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2230__A2 _1996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2014__A _2055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1974__D1 _1965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2518__B1 _2517_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3494__A1 _4132_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__B2 _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__B _4135_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output287_A _2860_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3706__C1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2859__A _2859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3681__C _3925_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2350_ _4250_/Q _3295_/C _2590_/B _2414_/A _3744_/B2 vssd1 vssd1 vccd1 vccd1 _2350_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2281_ _2380_/A vssd1 vssd1 vccd1 vccd1 _2281_/X sky130_fd_sc_hd__buf_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4020_ _4085_/CLK _4020_/D vssd1 vssd1 vccd1 vccd1 _4020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3788__A2 _2133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2460__A2 _2329_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1938__A _1938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4111__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1996_ _2018_/A vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__buf_2
X_3804_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3735_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4261__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3796_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2769__A _3489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2617_ _2380_/X _2614_/Y _2509_/A _2615_/Y _2616_/Y vssd1 vssd1 vccd1 vccd1 _2617_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _4191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2548_ _2542_/X _2547_/Y _2499_/X _2524_/X vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2920__A0 _4318_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4218_ _4262_/CLK _4218_/D vssd1 vssd1 vccd1 vccd1 _4218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ _3541_/B _2362_/X _2473_/Y _2478_/Y vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__3476__A1 _4124_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3476__B2 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2279__A2 _2245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4149_ _4389_/CLK _4149_/D vssd1 vssd1 vccd1 vccd1 _4149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3779__A2 _3764_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2451__A2 _2449_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2203__A2 _1961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2463__B1_N _4158_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__A2 _2260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2679__A _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2911__A0 _3250_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input46_A cpu_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3303__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4134__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output202_A _2976_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3957__B _3973_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2442__A2 _2438_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4284__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3520_ _3547_/A vssd1 vssd1 vccd1 vccd1 _3549_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3973__A _3973_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1953__A1 _1952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3155__A0 _3174_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2589__A _4275_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3451_ _3451_/A _3459_/B _3455_/C vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__and3_1
X_2402_ _3730_/A _2428_/A _2429_/A _2434_/A _4390_/Q vssd1 vssd1 vccd1 vccd1 _2402_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3382_ _3382_/A vssd1 vssd1 vccd1 vccd1 _4087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2333_ _2256_/X _2258_/X _2311_/X _2260_/X _4362_/Q vssd1 vssd1 vccd1 vccd1 _2333_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2264_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2453_/A sky130_fd_sc_hd__clkbuf_4
X_2195_ _4250_/Q vssd1 vssd1 vccd1 vccd1 _3023_/A sky130_fd_sc_hd__buf_2
XFILLER_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4003_/A vssd1 vssd1 vccd1 vccd1 _4388_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3213__A _3221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2969__B1 _3664_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2433__A2 _2432_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3867__B _3877_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3586__C _3586_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3883__A _3883_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1979_ input4/X vssd1 vssd1 vccd1 vccd1 _1983_/A sky130_fd_sc_hd__inv_2
XFILLER_101_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3718_ _3718_/A vssd1 vssd1 vccd1 vccd1 _4245_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3933__A2 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3649_ _3649_/A vssd1 vssd1 vccd1 vccd1 _4213_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2499__A _2499_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4007__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4157__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3123__A _3123_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2672__A2 _2133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input100_A gpio_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3496__C _3502_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4104__D _4104_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3793__A _3793_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__A2 _3902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3017__B _4240_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3688__B2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3688__A1 _4230_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2360__A1 _2330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output152_A _2537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2648__C1 _2647_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3033__A _3033_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2575__C _2638_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__A _3991_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2872__A _2888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2951_ _3174_/B _4078_/Q _3161_/A vssd1 vssd1 vccd1 vccd1 _3358_/C sky130_fd_sc_hd__mux2_4
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2882_ _3239_/C _4101_/Q _2916_/S vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__mux2_4
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4014__D _4014_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2179__A1 _1952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2811__S _2858_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3503_ _3503_/A vssd1 vssd1 vccd1 vccd1 _4137_/D sky130_fd_sc_hd__clkbuf_1
X_3434_ _3434_/A _3459_/B _3455_/C vssd1 vssd1 vccd1 vccd1 _3435_/A sky130_fd_sc_hd__and3_1
XANTENNA__2112__A _2129_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3128__A0 _3247_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3208__A _3221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__A1 _4226_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__B2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3365_ _3383_/A _3365_/B _3365_/C vssd1 vssd1 vccd1 vccd1 _3366_/A sky130_fd_sc_hd__or3_1
XANTENNA__2351__A1 _2343_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1951__A _1951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2351__B2 _2406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2316_ _2262_/X _2375_/A _2408_/A _2409_/A _2315_/Y vssd1 vssd1 vccd1 vccd1 _2316_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3296_ _2145_/C _2145_/D _3346_/C vssd1 vssd1 vccd1 vccd1 _4053_/D sky130_fd_sc_hd__a21oi_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2247_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3878__A _3878_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2178_ _4067_/Q _2093_/X _2177_/Y vssd1 vssd1 vccd1 vccd1 _2186_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2782__A _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3906__A2 _3902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3118__A _3118_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2022__A _2022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput102 gpio_dat_i[6] vssd1 vssd1 vccd1 vccd1 _2368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput113 spi_dat_i[13] vssd1 vssd1 vccd1 vccd1 _2483_/C sky130_fd_sc_hd__clkbuf_2
Xinput135 spi_dat_i[4] vssd1 vssd1 vccd1 vccd1 _2332_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput124 spi_dat_i[23] vssd1 vssd1 vccd1 vccd1 _2583_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2645__A2 _4178_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3938__D _3938_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3028__A _3032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4322__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2867__A _2867_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3150_ _3267_/B _4216_/Q _3150_/S vssd1 vssd1 vccd1 vccd1 _3655_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2333__A1 _2256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2333__B2 _2260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3081_ _3081_/A _3089_/B _3607_/C vssd1 vssd1 vccd1 vccd1 _3082_/A sky130_fd_sc_hd__and3_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2101_ _2237_/A vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__buf_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2032_ _4066_/Q vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2636__A2 _2428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2097__B1 _1962_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4009__D _4009_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3983_ _3983_/A vssd1 vssd1 vccd1 vccd1 _4374_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3210__B _3210_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2934_ _2934_/A vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__clkbuf_1
X_2865_ _3231_/B _4098_/Q _2911_/S vssd1 vssd1 vccd1 vccd1 _3407_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2232__B1_N _4179_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2796_ _2958_/S vssd1 vssd1 vccd1 vccd1 _2845_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2572__A1 _2572_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3417_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3437_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2777__A _2898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3348_ _4075_/Q _3314_/A _2063_/Y _3315_/A vssd1 vssd1 vccd1 vccd1 _4075_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3279_ _3328_/B _3279_/B _3279_/C _3286_/D vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__and4_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2627__A2 _2582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2943__C _3442_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3401__A _3401_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4001__A1 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4345__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2563__A1 _2419_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__B1 _2493_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3512__B1 _2767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2315__A1 _2313_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2618__A2 _2582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2079__B1 _2078_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3949__C _3963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3311__A _3311_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3030__B _4246_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2896_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2003__B1 _2002_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2554__A1 _2281_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2581_ _2581_/A vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3751__B1 _3735_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2554__B2 _2551_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4320_ _4391_/CLK _4320_/D vssd1 vssd1 vccd1 vccd1 _4320_/Q sky130_fd_sc_hd__dfxtp_1
X_4251_ _4251_/CLK _4251_/D vssd1 vssd1 vccd1 vccd1 _4251_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2306__B2 _2299_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2306__A1 _2281_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3202_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ _4250_/CLK _4182_/D vssd1 vssd1 vccd1 vccd1 _4182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3133_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3133_/X sky130_fd_sc_hd__clkbuf_1
X_3064_ _3064_/A vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4218__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2609__A2 _2366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2015_ _2055_/B vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3221__A _3221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2490__B1 _2404_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4368__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3966_ _3945_/D _3736_/Y _2255_/X _3724_/C _3992_/A vssd1 vssd1 vccd1 vccd1 _3966_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2917_ _2917_/A _2928_/B _3429_/A vssd1 vssd1 vccd1 vccd1 _2918_/A sky130_fd_sc_hd__and3_1
XANTENNA__2242__B1 _2346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3594__C _3594_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3897_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3942_/B sky130_fd_sc_hd__clkbuf_2
X_2848_ _2848_/A vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2545__A1 _2545_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2779_ _3190_/B _4084_/Q _2937_/S vssd1 vssd1 vccd1 vccd1 _3374_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4202__D _4202_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3891__A _3895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3742__B1 _3735_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2938__C _3439_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2300__A _2452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2233__B1 _2232_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__B1 _2510_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2784__A1 input61/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input76_A gpio_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__A1 _2526_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4112__D _4112_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__B2 _2534_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3733__B1 _2276_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3306__A _3953_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2210__A _2210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_10_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output232_A _3149_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3041__A _3041_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2583__C _2583_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2472__B1 _2471_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3976__A _3976_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3820_ _3820_/A vssd1 vssd1 vccd1 vccd1 _4298_/D sky130_fd_sc_hd__clkbuf_1
X_3751_ _4260_/Q _3750_/X _3735_/X _2440_/D _3738_/X vssd1 vssd1 vccd1 vccd1 _4260_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2702_ _2704_/A _4122_/Q vssd1 vssd1 vccd1 vccd1 _2703_/A sky130_fd_sc_hd__and2_1
X_3682_ _3682_/A vssd1 vssd1 vccd1 vccd1 _4227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2633_ _2328_/A _2329_/A _2469_/A _2632_/Y vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__o211a_1
Xoutput203 _2980_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[5] sky130_fd_sc_hd__buf_2
Xoutput225 _3130_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput214 _3094_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2527__A1 _2700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2564_ _2559_/X _2563_/Y _2499_/X _2524_/X vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4022__D _4022_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput247 _2658_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput258 _2668_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput236 _3061_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[5] sky130_fd_sc_hd__buf_2
X_4303_ _4346_/CLK _4303_/D vssd1 vssd1 vccd1 vccd1 _4303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput269 _2672_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[2] sky130_fd_sc_hd__buf_2
X_2495_ _2386_/X _2424_/X _4161_/Q vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3216__A _3216_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4234_ _4264_/CLK _4234_/D vssd1 vssd1 vccd1 vccd1 _4234_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4040__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2120__A _2120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4165_ _4177_/CLK _4165_/D vssd1 vssd1 vccd1 vccd1 _4165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _3241_/B _4206_/Q _3144_/S vssd1 vssd1 vccd1 vccd1 _3631_/C sky130_fd_sc_hd__mux2_1
XFILLER_83_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4180_/CLK _4096_/D vssd1 vssd1 vccd1 vccd1 _4096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4190__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3047_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3076_/S sky130_fd_sc_hd__buf_2
XANTENNA__3589__C _3600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3886__A _3886_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2766__A1 _4082_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3949_ _3949_/A _3973_/B _3963_/C vssd1 vssd1 vccd1 vccd1 _3950_/A sky130_fd_sc_hd__and3_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2230__A3 _3879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1974__C1 _1973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2518__A1 _2363_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2518__B2 _2450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3126__A _3126_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3479__C1 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2030__A _2030_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2965__A _3120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3494__A2 _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input130_A spi_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__C _3502_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4107__D _4107_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2904__S _2904_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3796__A _3796_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2206__B1 _2205_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output182_A _3003_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3706__B1 _3696_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2859__B _2872_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4063__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3036__A _3036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3681__D _3689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2280_ _2418_/A vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__buf_2
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3338__A_N _2158_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2693__A0 _3895_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4017__D _4017_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3803_ _3803_/A vssd1 vssd1 vccd1 vccd1 _4291_/D sky130_fd_sc_hd__clkbuf_1
X_1995_ _1951_/A _1994_/X _1942_/B vssd1 vssd1 vccd1 vccd1 _2018_/A sky130_fd_sc_hd__o21a_1
X_3734_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2115__A _4284_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3665_ _3665_/A vssd1 vssd1 vccd1 vccd1 _4220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2616_ _2407_/A _2406_/A _2324_/X _2552_/X _4385_/Q vssd1 vssd1 vccd1 vccd1 _2616_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__1954__A input6/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3596_ _3596_/A _3609_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__and3_1
X_2547_ _2419_/X _3550_/B _2546_/Y vssd1 vssd1 vccd1 vccd1 _2547_/Y sky130_fd_sc_hd__o21ai_1
X_2478_ _2474_/X _2452_/X _2453_/X _2454_/X _2477_/Y vssd1 vssd1 vccd1 vccd1 _2478_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__2920__A1 input54/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _4284_/CLK _4217_/D vssd1 vssd1 vccd1 vccd1 _4217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3476__A2 _3350_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2684__A0 _3283_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4148_ _4389_/CLK _4148_/D vssd1 vssd1 vccd1 vccd1 _4148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4251_/CLK _4079_/D vssd1 vssd1 vccd1 vccd1 _4079_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3779__A3 _3765_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2203__A3 _1918_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4086__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1947__C1 _1977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2911__A1 _4106_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input39_A cpu_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2385__A_N _2382_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__A0 _3279_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3303__B _3303_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3957__C _3963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3927__B1 _4346_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3973__B _3973_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1953__A2 _1932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _3450_/A vssd1 vssd1 vccd1 vccd1 _4114_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3155__A1 _4182_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3959__B1_N _2326_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2401_ _2450_/A vssd1 vssd1 vccd1 vccd1 _2434_/A sky130_fd_sc_hd__clkbuf_4
X_3381_ _3381_/A _3381_/B _3400_/C vssd1 vssd1 vccd1 vccd1 _3382_/A sky130_fd_sc_hd__and3_1
X_2332_ _2332_/A1 _2090_/A _2308_/X _2421_/A _2331_/Y vssd1 vssd1 vccd1 vccd1 _3530_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__4300__D _4300_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4002_ _4002_/A _4002_/B _4002_/C vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__and3_1
X_2263_ _2346_/A vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2809__S _2845_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2194_ _2128_/X _2133_/X _2780_/B vssd1 vssd1 vccd1 vccd1 _2194_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3213__B _3227_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2969__A1 _2197_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1949__A _4057_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3867__C _3867_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3717_ _3717_/A _4245_/Q _3721_/C _3724_/D vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__and4_1
X_1978_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2182_/B sky130_fd_sc_hd__buf_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3648_ _3648_/A _3661_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__and3_1
X_3579_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3600_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__4210__D _4210_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3404__A _3444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2657__A0 _3271_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3688__A2 _3351_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4120__D _4120_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2360__A2 _2424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4101__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3314__A _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output145_A _2460_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2648__B1 _2509_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output312_A _2948_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2575__D _2575_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2872__B _2872_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4251__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3073__A0 _3210_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2950_ _3794_/C _4008_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__mux2_2
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2881_ _3850_/A _4031_/Q _2905_/S vssd1 vssd1 vccd1 vccd1 _3239_/C sky130_fd_sc_hd__mux2_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2820__A0 _4301_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2179__A2 _1932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3502_ _3510_/A _4137_/Q _3502_/C vssd1 vssd1 vccd1 vccd1 _3503_/A sky130_fd_sc_hd__and3_1
XANTENNA__2112__B _2112_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3433_ _3433_/A vssd1 vssd1 vccd1 vccd1 _3459_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3128__A1 _4209_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3208__B _3227_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__A2 _3351_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4030__D _4030_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3383_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2887__A0 _3241_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2351__A2 _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2315_ _2313_/Y _2539_/A _2314_/Y vssd1 vssd1 vccd1 vccd1 _2315_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3224__A _3224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3295_ _3591_/A _3298_/A _3295_/C vssd1 vssd1 vccd1 vccd1 _3346_/C sky130_fd_sc_hd__or3_4
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2639__B1 _2638_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2246_ _2579_/A vssd1 vssd1 vccd1 vccd1 _2246_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _2038_/A _3902_/A _2176_/Y _1973_/X _2136_/X vssd1 vssd1 vccd1 vccd1 _2177_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2811__A0 _3208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4205__D _4205_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3894__A _3894_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2303__A _2429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4124__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2327__C1 _2125_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput103 gpio_dat_i[7] vssd1 vssd1 vccd1 vccd1 _2396_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput125 spi_dat_i[24] vssd1 vssd1 vccd1 vccd1 _2594_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput114 spi_dat_i[14] vssd1 vssd1 vccd1 vccd1 _2496_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput136 spi_dat_i[5] vssd1 vssd1 vccd1 vccd1 _2352_/D1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4274__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2973__A _3343_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2802__A0 _4298_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4115__D _4115_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3309__A _3309_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3028__B _4245_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output262_A _2736_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2318__C1 _2125_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2869__A0 _3845_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2333__A2 _2258_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3044__A _3044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2100_ _2106_/A _2112_/B _2099_/Y vssd1 vssd1 vccd1 vccd1 _2237_/A sky130_fd_sc_hd__o21ai_4
X_3080_ _3215_/B _4196_/Q _3109_/S vssd1 vssd1 vccd1 vccd1 _3607_/C sky130_fd_sc_hd__mux2_1
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2031_ _2031_/A _3320_/B _2031_/C vssd1 vssd1 vccd1 vccd1 _2085_/A sky130_fd_sc_hd__nor3_1
XANTENNA__2883__A _2888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2097__A1 _1949_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3982_ _3982_/A _3999_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__and3_1
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2933_ _2943_/A _3447_/B _3437_/C vssd1 vssd1 vccd1 vccd1 _2934_/A sky130_fd_sc_hd__and3_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3210__C _3224_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2822__S _2858_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4025__D _4025_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2864_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2911_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2795_ _4297_/Q input63/X _2844_/S vssd1 vssd1 vccd1 vccd1 _3817_/A sky130_fd_sc_hd__mux2_8
XANTENNA__4147__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3219__A _3224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2572__A2 _2444_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1962__A _1962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3416_ _3416_/A vssd1 vssd1 vccd1 vccd1 _4101_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4297__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3347_ _3347_/A vssd1 vssd1 vccd1 vccd1 _4074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3278_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3889__A _3889_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2793__A _2793_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2229_ _4180_/Q _2543_/A _2356_/C vssd1 vssd1 vccd1 vccd1 _2418_/A sky130_fd_sc_hd__o21ai_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3129__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4001__A2 _3992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2548__C1 _2524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3760__A1 _3752_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2563__A2 _3552_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3512__A1 _4142_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3512__B2 _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2315__A2 _2539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input21_A cpu_adr_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__A _3799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2079__A1 _4349_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2208__A _2208_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2003__A1 input33/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2554__A2 _2550_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2580_ _2512_/X _2513_/X _3989_/A _2579_/X vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3751__A1 _4260_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2878__A _2888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__B2 _2440_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4250_ _4250_/CLK _4250_/D vssd1 vssd1 vccd1 vccd1 _4250_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2306__A2 _2291_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4181_ _4251_/CLK _4181_/D vssd1 vssd1 vccd1 vccd1 _4181_/Q sky130_fd_sc_hd__dfxtp_1
X_3201_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3297_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3132_ _3135_/A _3142_/B _3642_/C vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__and3_1
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3063_ _3063_/A _3070_/B _3596_/A vssd1 vssd1 vccd1 vccd1 _3064_/A sky130_fd_sc_hd__and3_1
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2817__S _2851_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3502__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2014_ _2055_/A vssd1 vssd1 vccd1 vccd1 _2136_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3221__B _3227_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2490__A1 _2482_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3965_ _3965_/A vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1957__A _2022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2242__B2 _2257_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2242__A1 _2117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2916_ _3253_/C _4107_/Q _2916_/S vssd1 vssd1 vccd1 vccd1 _3429_/A sky130_fd_sc_hd__mux2_2
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3896_ _3896_/A vssd1 vssd1 vccd1 vccd1 _4330_/D sky130_fd_sc_hd__clkbuf_1
X_2847_ _2859_/A _2872_/B _3400_/A vssd1 vssd1 vccd1 vccd1 _2848_/A sky130_fd_sc_hd__and3_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2778_ _3810_/C _4014_/Q _2826_/S vssd1 vssd1 vccd1 vccd1 _3190_/B sky130_fd_sc_hd__mux2_2
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3891__B _3935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2788__A _2788_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2545__A2 _3369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3742__B2 input99/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3742__A1 _4254_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4389_/CLK _4379_/D vssd1 vssd1 vccd1 vccd1 _4379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3412__A _3461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4312__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2028__A _2028_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2233__A1 _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3981__A1 _4373_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2536__A2 _2532_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3733__A1 _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input69_A cpu_sel_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2210__B _2210_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output225_A _3130_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__A1 _2472_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2209__D1 _3301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3750_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2701_ _2739_/A vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ _3699_/A _4227_/Q _3925_/D _3689_/D vssd1 vssd1 vccd1 vccd1 _3682_/A sky130_fd_sc_hd__and4_1
XANTENNA__3992__A _3992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4303__D _4303_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2632_ _2526_/X _2629_/Y _2509_/X _2630_/Y _2631_/Y vssd1 vssd1 vccd1 vccd1 _2632_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput226 _3133_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput215 _3097_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput204 _2982_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__2527__A2 _2678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2563_ _2419_/X _3552_/B _2562_/Y vssd1 vssd1 vccd1 vccd1 _2563_/Y sky130_fd_sc_hd__o21ai_1
Xoutput259 _2730_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput248 _2708_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput237 _3064_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__2401__A _2450_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4302_ _4302_/CLK _4302_/D vssd1 vssd1 vccd1 vccd1 _4302_/Q sky130_fd_sc_hd__dfxtp_1
X_4233_ _4264_/CLK _4233_/D vssd1 vssd1 vccd1 vccd1 _4233_/Q sky130_fd_sc_hd__dfxtp_1
X_2494_ _2406_/X _2407_/X _2408_/X _2409_/X _2493_/Y vssd1 vssd1 vccd1 vccd1 _2494_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _4177_/CLK _4164_/D vssd1 vssd1 vccd1 vccd1 _4164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3115_ _3115_/A vssd1 vssd1 vccd1 vccd1 _3144_/S sky130_fd_sc_hd__buf_2
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4095_ _4199_/CLK _4095_/D vssd1 vssd1 vccd1 vccd1 _4095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3063_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3232__A _3232_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4335__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2463__A1 _2287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3948_ _4002_/C vssd1 vssd1 vccd1 vccd1 _3963_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4213__D _4213_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3879_ _3879_/A _3893_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__and3_1
XANTENNA__1974__B1 _1971_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2518__A2 _2449_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3407__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2311__A _2517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3479__B1 _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2030__B _2030_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2151__B1 _4351_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3142__A _3151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input123_A spi_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__B _3796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2206__A1 _2662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4123__D _4123_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2920__S _2940_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3706__A1 _4238_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3706__B2 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4208__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2859__C _3405_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2221__A _2450_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3317__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output175_A _2443_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3036__B _4249_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4358__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2142__B1 _4335_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3052__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2693__A1 _4050_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3802_ _3802_/A _3821_/B _3903_/A vssd1 vssd1 vccd1 vccd1 _3803_/A sky130_fd_sc_hd__and3_1
X_1994_ _1994_/A vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__buf_2
X_3733_ _3727_/X _3729_/X _3732_/X _2276_/Y _3566_/X vssd1 vssd1 vccd1 vccd1 _4251_/D
+ sky130_fd_sc_hd__o311a_1
X_3664_ _3798_/A _3673_/B _3664_/C vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__or3_1
XANTENNA__4033__D _4033_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2615_ _4278_/Q _2322_/X _2298_/A input93/X vssd1 vssd1 vccd1 vccd1 _2615_/Y sky130_fd_sc_hd__a22oi_4
X_3595_ _3595_/A vssd1 vssd1 vccd1 vccd1 _4190_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2131__A _2678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3227__A _3247_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2546_ _2427_/X _2428_/X _2303_/X _2304_/X _4376_/Q vssd1 vssd1 vccd1 vccd1 _2546_/Y
+ sky130_fd_sc_hd__o221ai_1
X_4393__319 vssd1 vssd1 vccd1 vccd1 _4393__319/HI cpu_rty_o sky130_fd_sc_hd__conb_1
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2477_ _2475_/Y _2366_/X _2476_/Y vssd1 vssd1 vccd1 vccd1 _2477_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__1970__A _1970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4216_ _4264_/CLK _4216_/D vssd1 vssd1 vccd1 vccd1 _4216_/Q sky130_fd_sc_hd__dfxtp_1
X_4147_ _4389_/CLK _4147_/D vssd1 vssd1 vccd1 vccd1 _4147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2684__A1 _4118_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4250_/CLK _4078_/D vssd1 vssd1 vccd1 vccd1 _4078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3897__A _3897_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3029_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4208__D _4208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1947__B1 _1946_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3137__A _3137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__A1 _4117_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3303__C _3317_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4118__D _4118_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2915__S _2936_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3600__A _3600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2216__A _3127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output292_A _2884_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4030__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3927__A1 _2121_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3973__C _3996_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4180__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2400_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2428_/A sky130_fd_sc_hd__buf_4
XANTENNA__3047__A _3120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3380_ _3444_/A vssd1 vssd1 vccd1 vccd1 _3400_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2331_ _2330_/X _2424_/A _4151_/Q vssd1 vssd1 vccd1 vccd1 _2331_/Y sky130_fd_sc_hd__a21boi_1
X_2262_ _3730_/B vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__buf_4
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4001_ _3991_/X _3992_/X _2632_/Y vssd1 vssd1 vccd1 vccd1 _4387_/D sky130_fd_sc_hd__o21bai_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2193_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2780_/B sky130_fd_sc_hd__buf_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3213__C _3213_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4028__D _4028_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2825__S _2825_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3510__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2969__A2 _2200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2126__A _4146_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3716_ _4244_/Q _3167_/B _3044_/A _3697_/A _3705_/X vssd1 vssd1 vccd1 vccd1 _4244_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1965__A _2055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1977_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3647_ _3647_/A vssd1 vssd1 vccd1 vccd1 _4212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3578_ _3578_/A vssd1 vssd1 vccd1 vccd1 _3680_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3551__C1 _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2529_ _2529_/A vssd1 vssd1 vccd1 vccd1 _2628_/A sky130_fd_sc_hd__buf_2
XANTENNA__2796__A _2958_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2657__A1 _4114_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3420__A _3420_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4053__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2036__A _4067_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3542__C1 _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input51_A cpu_dat_i[24] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2648__B2 _2646_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2648__A1 _2526_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2872__C _3410_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output305_A _2781_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3330__A _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3073__A1 _4194_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2880_ _4311_/Q input47/X _2904_/S vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__mux2_8
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2820__A1 input36/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2584__B1 _2583_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3501_ _4136_/Q _3488_/X _3489_/X _3490_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _4136_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3781__C1 _3774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3432_ _3432_/A vssd1 vssd1 vccd1 vccd1 _4108_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4311__D _4311_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3208__C _3208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3533__C1 _3562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3363_ _3591_/A vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2887__A1 _4102_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2314_ _2412_/A _2590_/B _2414_/A _2314_/D vssd1 vssd1 vccd1 vccd1 _2314_/Y sky130_fd_sc_hd__nand4_2
X_3294_ _3315_/A _3294_/B _3294_/C vssd1 vssd1 vccd1 vccd1 _4052_/D sky130_fd_sc_hd__nand3_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2639__A1 _2637_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2245_ _2329_/A vssd1 vssd1 vccd1 vccd1 _2245_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3224__B _3224_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4076__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2176_ _2121_/A _2160_/X _4347_/Q vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3240__A _3240_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2811__A1 _4089_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4221__D _4221_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2327__B1 _2326_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3415__A _3415_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput126 spi_dat_i[25] vssd1 vssd1 vccd1 vccd1 _3557_/A1 sky130_fd_sc_hd__buf_2
Xinput115 spi_dat_i[15] vssd1 vssd1 vccd1 vccd1 _2503_/C sky130_fd_sc_hd__clkbuf_2
Xinput104 gpio_dat_i[8] vssd1 vssd1 vccd1 vccd1 _2415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput137 spi_dat_i[6] vssd1 vssd1 vccd1 vccd1 _2361_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2802__A1 input64/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input99_A gpio_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2566__B1 _2565_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__C1 _3755_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4131__D _4131_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3515__C1 _3504_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2318__B1 _3957_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output255_A _2723_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2869__A1 _4029_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4099__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3044__B _3052_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2030_ _2030_/A _2030_/B _2030_/C _2030_/D vssd1 vssd1 vccd1 vccd1 _2031_/C sky130_fd_sc_hd__nand4_1
XANTENNA__2883__B _2901_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2097__A2 _2093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3060__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3981_ _4373_/Q _3965_/X _2510_/Y _3966_/Y vssd1 vssd1 vccd1 vccd1 _4373_/D sky130_fd_sc_hd__a211o_1
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2932_ _3262_/B _4110_/Q _2942_/S vssd1 vssd1 vccd1 vccd1 _3437_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4306__D _4306_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3210__D _3219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2863_ _3843_/C _4028_/Q _2886_/S vssd1 vssd1 vccd1 vccd1 _3231_/B sky130_fd_sc_hd__mux2_4
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2404__A _2499_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2794_ _2957_/S vssd1 vssd1 vccd1 vccd1 _2844_/S sky130_fd_sc_hd__buf_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3219__B _3219_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2572__A3 _2514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4041__D _4041_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1962__B _1962_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4395_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3415_ _3415_/A _3429_/B _3424_/C vssd1 vssd1 vccd1 vccd1 _3416_/A sky130_fd_sc_hd__and3_1
XANTENNA__3235__A _3235_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3346_ _3346_/A _3346_/B _3346_/C vssd1 vssd1 vccd1 vccd1 _3347_/A sky130_fd_sc_hd__or3_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3277_ _3277_/A vssd1 vssd1 vccd1 vccd1 _4046_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3889__B _3893_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2228_ _4285_/Q _2130_/A _3945_/D vssd1 vssd1 vccd1 vccd1 _2356_/C sky130_fd_sc_hd__o21a_1
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2159_ _2159_/A _2159_/B vssd1 vssd1 vccd1 vccd1 _2211_/A sky130_fd_sc_hd__nor2_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4216__D _4216_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2314__A _2412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3129__B _3142_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3745__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2548__B1 _2499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4241__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3145__A _3151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3512__A2 _3308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4391__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2079__A2 _2012_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A cpu_adr_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4126__D _4126_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2224__A _2328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2003__A2 _2001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__A2 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2878__B _2901_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3055__A _3657_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4180_ _4180_/CLK _4180_/D vssd1 vssd1 vccd1 vccd1 _4180_/Q sky130_fd_sc_hd__dfxtp_2
X_3200_ _3200_/A vssd1 vssd1 vccd1 vccd1 _4017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3131_ _3250_/B _4210_/Q _3144_/S vssd1 vssd1 vccd1 vccd1 _3642_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2894__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3062_ _3199_/C _4191_/Q _3076_/S vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3502__B _4137_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2013_ _1930_/X _1932_/X _4342_/Q vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_63_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3221__C _3221_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2490__A2 _2489_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2833__S _2858_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4036__D _4036_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4114__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3964_ _3964_/A vssd1 vssd1 vccd1 vccd1 _4364_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2778__A0 _3810_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2242__A2 _2344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__C1 _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2915_ _3865_/A _4037_/Q _2936_/S vssd1 vssd1 vccd1 vccd1 _3253_/C sky130_fd_sc_hd__mux2_2
X_3895_ _3895_/A _3935_/B _3895_/C vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__or3_1
X_2846_ _3221_/C _4095_/Q _2858_/S vssd1 vssd1 vccd1 vccd1 _3400_/A sky130_fd_sc_hd__mux2_4
XANTENNA__2134__A _2134_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1986__D1 _1985_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4264__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2777_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2826_/S sky130_fd_sc_hd__buf_2
XANTENNA__1973__A _2055_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2545__A3 _2286_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3742__A2 _3734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2950__A0 _3794_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3891__C _3891_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _4390_/CLK _4378_/D vssd1 vssd1 vccd1 vccd1 _4378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input6_A cpu_adr_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3329_/A vssd1 vssd1 vccd1 vccd1 _4067_/D sky130_fd_sc_hd__clkbuf_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2028__B _2072_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2233__A2 _2190_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__A2 _3965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2044__A _2044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3733__A2 _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2941__A0 _3877_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3603__A _3603_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4137__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2219__A _2257_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output218_A _3107_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2472__A2 _2444_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2209__C1 _1990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4287__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2700_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2739_/A sky130_fd_sc_hd__clkbuf_4
X_3680_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2889__A _2889_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2631_ _2481_/X _2501_/X _2429_/X _2430_/X _4387_/Q vssd1 vssd1 vccd1 vccd1 _2631_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput205 _2984_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[7] sky130_fd_sc_hd__buf_2
Xoutput216 _3100_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2436__A_N _2382_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2562_ _2427_/X _2428_/X _2303_/X _2304_/X _4378_/Q vssd1 vssd1 vccd1 vccd1 _2562_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput227 _3136_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput238 _3068_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput249 _2710_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[11] sky130_fd_sc_hd__buf_2
XANTENNA__2932__A0 _3262_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4301_ _4346_/CLK _4301_/D vssd1 vssd1 vccd1 vccd1 _4301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _4264_/CLK _4232_/D vssd1 vssd1 vccd1 vccd1 _4232_/Q sky130_fd_sc_hd__dfxtp_1
X_2493_ _2491_/Y _2411_/X _2492_/Y vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3513__A _3516_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4163_ _4180_/CLK _4163_/D vssd1 vssd1 vccd1 vccd1 _4163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3114_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3114_/X sky130_fd_sc_hd__clkbuf_1
X_4094_ _4180_/CLK _4094_/D vssd1 vssd1 vccd1 vccd1 _4094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3045_ _3045_/A vssd1 vssd1 vccd1 vccd1 _3045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2129__A _2129_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2463__A2 _3468_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1968__A _4056_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3947_ _3976_/A vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ _3878_/A vssd1 vssd1 vccd1 vccd1 _4322_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1974__A1 _4336_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2829_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2799__A _2799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3407__B _3413_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3479__A1 _4126_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3479__B2 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2030__C _2030_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3423__A _3423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2151__A1 _2121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3142__B _3142_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2039__A _2059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input116_A spi_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__C _3903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2206__A2 _3914_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input81_A gpio_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2611__C1 _2610_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3706__A2 _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2914__A0 _4317_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3317__B _3317_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output168_A _2649_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2142__A1 _2121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3052__B _3052_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3801_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3821_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4314__D _4314_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _2204_/A vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2602__C1 _2601_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3732_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3732_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3663_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3798_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3158__B1 _3574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3508__A _3508_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2614_ _3559_/A1 _2420_/X _2421_/X _2613_/Y vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__2412__A _2412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3594_ _3611_/A _3611_/B _3594_/C vssd1 vssd1 vccd1 vccd1 _3595_/A sky130_fd_sc_hd__or3_1
XANTENNA__2905__A0 _3861_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3227__B _3227_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2545_ _2545_/A1 _3369_/A _2286_/A _2544_/Y vssd1 vssd1 vccd1 vccd1 _3550_/B sky130_fd_sc_hd__a31oi_4
XFILLER_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4302__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2476_ _2575_/A _2520_/B _2520_/C _2476_/D vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__nand4_2
X_4215_ _4275_/CLK _4215_/D vssd1 vssd1 vccd1 vccd1 _4215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _4177_/CLK _4146_/D vssd1 vssd1 vccd1 vccd1 _4146_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3243__A _3247_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4251_/CLK _4077_/D vssd1 vssd1 vccd1 vccd1 _4077_/Q sky130_fd_sc_hd__dfxtp_1
X_3028_ _3032_/A _4245_/Q vssd1 vssd1 vccd1 vccd1 _3029_/A sky130_fd_sc_hd__and2_1
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4224__D _4224_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1947__A1 _1939_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3418__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2322__A _3720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2992__A _2992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3303__D _3326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3600__B _3609_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4134__D _4134_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2931__S _2941_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3927__A2 _2201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2060__B1 _2059_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output285_A _2848_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4325__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3328__A _3328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__buf_2
X_2261_ _2256_/X _2258_/X _3728_/A _2260_/X _4358_/Q vssd1 vssd1 vccd1 vccd1 _2261_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_69_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3063__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _4386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2192_ _2782_/A vssd1 vssd1 vccd1 vccd1 _2903_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4309__D _4309_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3213__D _3234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3510__B _4141_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2407__A _2407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4044__D _4044_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1976_ _4055_/Q vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__inv_2
X_3715_ _3715_/A vssd1 vssd1 vccd1 vccd1 _4243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3238__A _3264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3646_ _3659_/A _3659_/B _3646_/C vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__or3_1
XANTENNA__2339__D1 _2338_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _4184_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1981__A _2078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3551__B1 _2549_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2528_ _3428_/A vssd1 vssd1 vccd1 vccd1 _3466_/C sky130_fd_sc_hd__clkbuf_4
X_2459_ _3539_/B _2362_/X _2451_/Y _2458_/Y vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__o211ai_4
XFILLER_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4129_ _4177_/CLK _4129_/D vssd1 vssd1 vccd1 vccd1 _4129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4219__D _4219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3420__B _3429_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4348__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2042__B1 _4064_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3148__A _3151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2593__A1 _2386_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2987__A _2987_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3542__B1 _2484_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input44_A cpu_dat_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2648__A2 _2645_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4129__D _4129_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2926__S _2936_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3611__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output200_A _3037_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2661__S _2935_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3058__A _3058_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3500_ _3500_/A vssd1 vssd1 vccd1 vccd1 _4135_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2584__A1 _3466_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2584__B2 _3544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__B1 _2624_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3431_ _3431_/A _3437_/B _3431_/C vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__or3_1
XANTENNA__3208__D _3208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3533__B1 _2388_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3362_ _3362_/A vssd1 vssd1 vccd1 vccd1 _4079_/D sky130_fd_sc_hd__clkbuf_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2313_ _4253_/Q vssd1 vssd1 vccd1 vccd1 _2313_/Y sky130_fd_sc_hd__inv_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3293_ _3293_/A _3335_/A _3707_/A vssd1 vssd1 vccd1 vccd1 _3315_/A sky130_fd_sc_hd__and3_2
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2639__A2 _2366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2244_ _2582_/A vssd1 vssd1 vccd1 vccd1 _2329_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3224__C _3224_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4039__D _4039_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2175_ _2175_/A _2175_/B _2175_/C _3317_/B vssd1 vssd1 vccd1 vccd1 _2187_/A sky130_fd_sc_hd__nand4_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3521__A _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2137__A _2137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1976__A _4055_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1959_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__buf_2
X_3629_ _3629_/A _3633_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__and3_1
XANTENNA__2327__A1 _2224_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3415__B _3429_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput127 spi_dat_i[26] vssd1 vssd1 vccd1 vccd1 _2605_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput116 spi_dat_i[16] vssd1 vssd1 vccd1 vccd1 _2516_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput105 gpio_dat_i[9] vssd1 vssd1 vccd1 vccd1 _2440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput138 spi_dat_i[7] vssd1 vssd1 vccd1 vccd1 _2385_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__4020__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3431__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4170__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A1 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2566__A1 _3553_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__B1 _3754_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3515__B1 _2767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2318__A1 _2224_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3606__A _3606_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output248_A _2708_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output150_A _2511_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3044__C _3582_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2883__C _3415_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3060__B _3070_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3980_ _3968_/X _3969_/X _2494_/X _2498_/Y vssd1 vssd1 vccd1 vccd1 _4372_/D sky130_fd_sc_hd__o22a_1
XFILLER_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2254__B1 _2253_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2931_ _3871_/C _4040_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _3262_/B sky130_fd_sc_hd__mux2_4
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2862_ _4308_/Q input43/X _2885_/S vssd1 vssd1 vccd1 vccd1 _3843_/C sky130_fd_sc_hd__mux2_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2793_ _2793_/A vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4322__D _4322_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3219__C _3224_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3516__A _3516_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2420__A _3441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2572__A4 _2445_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2309__A1 _2644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3414_ _3414_/A vssd1 vssd1 vccd1 vccd1 _4100_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1962__C _1962_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4043__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _4073_/Q _3314_/A _2059_/Y _3315_/A vssd1 vssd1 vccd1 vccd1 _4073_/D sky130_fd_sc_hd__o211a_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3276_ _3276_/A _3276_/B _3276_/C _3317_/C vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__or4_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2225_/Y _2683_/A _2446_/A vssd1 vssd1 vccd1 vccd1 _2543_/A sky130_fd_sc_hd__a21boi_4
XFILLER_86_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3889__C _3914_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3251__A _3251_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4193__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2493__B1 _2492_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2158_ _2158_/A _2158_/B _2158_/C _2158_/D vssd1 vssd1 vccd1 vccd1 _2159_/B sky130_fd_sc_hd__nand4_1
X_2089_ _2529_/A vssd1 vssd1 vccd1 vccd1 _2090_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2314__B _2590_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3129__C _3638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4232__D _4232_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3745__B1 _2369_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2548__A1 _2542_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3426__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__A3 _3748_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2330__A _2422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3145__B _3657_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3161__A _3161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2236__B1 _2213_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4142__D _4142_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output198_A _2969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3736__B1 _2453_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4066__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2878__C _3413_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3336__A input1/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_13_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4250_/CLK sky130_fd_sc_hd__clkbuf_16
X_3130_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2894__B _2901_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3071__A _3071_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3061_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3502__C _3502_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2012_ _2167_/A _2012_/B vssd1 vssd1 vccd1 vccd1 _2012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4317__D _4317_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3221__D _3234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3963_ _3963_/A _3973_/B _3963_/C vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__and3_1
XANTENNA__2778__A1 _4014_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2415__A _2507_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__B1 _2468_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2914_ _4317_/Q input53/X _2935_/S vssd1 vssd1 vccd1 vccd1 _3865_/A sky130_fd_sc_hd__mux2_4
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _4329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2845_ _3837_/A _4025_/Q _2845_/S vssd1 vssd1 vccd1 vccd1 _3221_/C sky130_fd_sc_hd__mux2_2
XANTENNA__1986__C1 _2137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4052__D _4052_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2776_ _4294_/Q input60/X _2825_/S vssd1 vssd1 vccd1 vccd1 _3810_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3246__A _3246_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2150__A _2150_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2950__A1 _4008_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4377_ _4389_/CLK _4377_/D vssd1 vssd1 vccd1 vccd1 _4377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _3328_/A _3328_/B _3695_/A _3925_/D vssd1 vssd1 vccd1 vccd1 _3329_/A sky130_fd_sc_hd__and4_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _3692_/A vssd1 vssd1 vccd1 vccd1 _3279_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2598__B1_N _4172_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4227__D _4227_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2028__C _2081_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__A3 _2231_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3966__B1 _3992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4089__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2044__B _2081_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3733__A3 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2941__A1 _4042_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2995__A _2999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2457__B1 _2456_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4137__D _4137_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2472__A3 _2308_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2209__B1 _1974_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2235__A _2638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2630_ _4280_/Q _2295_/X _2298_/X input95/X vssd1 vssd1 vccd1 vccd1 _2630_/Y sky130_fd_sc_hd__a22oi_4
Xoutput217 _3104_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput206 _2987_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[8] sky130_fd_sc_hd__buf_2
X_2561_ _2561_/A1 _3369_/A _2286_/A _2560_/Y vssd1 vssd1 vccd1 vccd1 _3552_/B sky130_fd_sc_hd__a31oi_4
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput228 _3140_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput239 _3071_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[8] sky130_fd_sc_hd__buf_2
XANTENNA__2932__A1 _4110_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2492_ _2590_/A _2557_/B _2590_/C _2492_/D vssd1 vssd1 vccd1 vccd1 _2492_/Y sky130_fd_sc_hd__nand4_2
XANTENNA_clkbuf_leaf_20_CLK_A _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _4326_/CLK _4300_/D vssd1 vssd1 vccd1 vccd1 _4300_/Q sky130_fd_sc_hd__dfxtp_1
X_4231_ _4264_/CLK _4231_/D vssd1 vssd1 vccd1 vccd1 _4231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4162_ _4172_/CLK _4162_/D vssd1 vssd1 vccd1 vccd1 _4162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2696__A0 _4331_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3513__B _4143_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3113_ _3117_/A _3125_/B _3629_/A vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__and3_1
X_4093_ _4225_/CLK _4093_/D vssd1 vssd1 vccd1 vccd1 _4093_/Q sky130_fd_sc_hd__dfxtp_1
X_3044_ _3044_/A _3052_/B _3582_/C vssd1 vssd1 vccd1 vccd1 _3045_/A sky130_fd_sc_hd__and3_1
XANTENNA__2448__B1 _2447_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2129__B _2129_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4047__D _4047_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2844__S _2844_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4231__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3946_ _3946_/A vssd1 vssd1 vccd1 vccd1 _4357_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2145__A _3294_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2620__B1 _2619_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3877_ _3895_/A _3877_/B _3877_/C vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__or3_1
XANTENNA__1984__A _2055_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1974__A2 _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2828_ _2828_/A _2841_/B _3394_/C vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__and3_1
XANTENNA__2799__B _2812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4381__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2759_ _3197_/A vssd1 vssd1 vccd1 vccd1 _2955_/S sky130_fd_sc_hd__buf_2
XANTENNA__3407__C _3407_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3479__A2 _3350_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3704__A _3704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2030__D _2030_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2687__A0 _4329_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2151__A2 _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3142__C _3648_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input109_A spi_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__B1 _2062_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2055__A _2055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2611__B1 _2606_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input74_A gpio_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2914__A1 input53/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3317__C _3317_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4104__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3614__A _3614_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output230_A _3146_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2142__A2 _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3052__C _3586_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4254__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2664__S _2936_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2850__A0 _3839_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _3800_/A vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _3765_/A vssd1 vssd1 vccd1 vccd1 _3748_/A sky130_fd_sc_hd__clkbuf_2
X_1992_ _4076_/Q vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2602__B1 _2293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3662_ _3662_/A vssd1 vssd1 vccd1 vccd1 _4219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3158__A1 _2988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2613_ _2319_/X _2248_/X _4174_/Q vssd1 vssd1 vccd1 vccd1 _2613_/Y sky130_fd_sc_hd__a21boi_1
X_3593_ _3617_/A vssd1 vssd1 vccd1 vccd1 _3611_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2544_ _2386_/X _2424_/X _4165_/Q vssd1 vssd1 vccd1 vccd1 _2544_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__2905__A1 _4035_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3227__C _3227_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4330__D _4330_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3524__A _3544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2475_ _4263_/Q vssd1 vssd1 vccd1 vccd1 _2475_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2839__S _2886_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4214_ _4282_/CLK _4214_/D vssd1 vssd1 vccd1 vccd1 _4214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2669__A0 _4326_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4145_ _4250_/CLK _4145_/D vssd1 vssd1 vccd1 vccd1 _4145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__B _3253_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4076_ _4391_/CLK _4076_/D vssd1 vssd1 vccd1 vccd1 _4076_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1979__A input4/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3027_ _3027_/A vssd1 vssd1 vccd1 vccd1 _3027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3929_ _4347_/Q _3908_/A _2038_/Y _3909_/X _3903_/X vssd1 vssd1 vccd1 vccd1 _4347_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__1947__A2 _2168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3418__B _3437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4127__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4240__D _4240_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3434__A _3434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4277__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3085__A0 _3217_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3600__C _3600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__A0 _3831_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__A3 _1994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2513__A _2582_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3609__A _3609_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2060__A1 _4073_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output180_A _2998_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3328__B _3328_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4150__D _4150_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output278_A _2705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2899__A0 _3858_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3344__A _3344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2260_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2260_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3063__B _3070_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2191_ _2139_/Y _2864_/A _2190_/Y vssd1 vssd1 vccd1 vccd1 _2782_/A sky130_fd_sc_hd__o21ai_1
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3076__A0 _3213_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3510__C _3657_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4325__D _4325_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1968_/Y _3332_/A _1974_/Y vssd1 vssd1 vccd1 vccd1 _3303_/B sky130_fd_sc_hd__o21ai_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3714_ _3717_/A _4243_/Q _3721_/C _3724_/D vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__and4_1
XANTENNA__2423__A _2423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__C1 _2586_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2339__C1 _2409_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3645_ _3645_/A vssd1 vssd1 vccd1 vccd1 _4211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4060__D _4060_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3576_ _3586_/A _3586_/B _3576_/C vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__or3_1
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3551__A1 _3551_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2527_ _2700_/A _2678_/A _2387_/A vssd1 vssd1 vccd1 vccd1 _3428_/A sky130_fd_sc_hd__o21ai_2
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2458_ _2262_/X _2452_/X _2453_/X _2454_/X _2457_/Y vssd1 vssd1 vccd1 vccd1 _2458_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__3254__A _3254_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2389_ _3536_/A _2385_/X _2388_/Y vssd1 vssd1 vccd1 vccd1 _2389_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2511__C1 _2469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _4177_/CLK _4128_/D vssd1 vssd1 vccd1 vccd1 _4128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4059_ _4326_/CLK _4059_/D vssd1 vssd1 vccd1 vccd1 _4059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3420__C _3424_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4235__D _4235_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2290__A1 _2287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2578__C1 _2577_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3429__A _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2042__A1 _1993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2593__A2 _2289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3148__B _3657_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3542__A1 _2483_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3164__A input1/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A cpu_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2502__C1 _4373_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3611__B _3611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2805__A0 _3204_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4145__D _4145_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2942__S _2942_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2569__C1 _2568_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3339__A _3339_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2033__A1 _2120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2584__A2 _4170_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__A1 _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3430_ _3430_/A vssd1 vssd1 vccd1 vccd1 _4107_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3533__A1 _2385_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3361_ _3361_/A _3381_/B _3376_/C vssd1 vssd1 vccd1 vccd1 _3362_/A sky130_fd_sc_hd__and3_1
XANTENNA__3074__A _3081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _2256_/X _2258_/X _2311_/X _2260_/X _4360_/Q vssd1 vssd1 vccd1 vccd1 _2312_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3292_ _3292_/A vssd1 vssd1 vccd1 vccd1 _4051_/D sky130_fd_sc_hd__clkbuf_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2418_/A _3564_/A _2239_/Y _2292_/A vssd1 vssd1 vccd1 vccd1 _2582_/A sky130_fd_sc_hd__o22ai_4
XANTENNA__3224__D _3245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3802__A _3802_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2174_ _2171_/Y _2153_/C _2173_/Y vssd1 vssd1 vccd1 vccd1 _3317_/B sky130_fd_sc_hd__o21ai_2
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2418__A _2418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4055__D _4055_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2009__D1 _1985_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3249__A _3343_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2153__A _2153_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1958_ _2078_/C vssd1 vssd1 vccd1 vccd1 _1971_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__1992__A _4076_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3628_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3648_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2327__A2 _2245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3559_ _3559_/A1 _3365_/B _3544_/X _2613_/Y _3547_/X vssd1 vssd1 vccd1 vccd1 _4174_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 gpio_err_i vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput117 spi_dat_i[17] vssd1 vssd1 vccd1 vccd1 _2530_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__3415__C _3424_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput128 spi_dat_i[27] vssd1 vssd1 vccd1 vccd1 _3559_/A1 sky130_fd_sc_hd__buf_2
Xinput139 spi_dat_i[8] vssd1 vssd1 vccd1 vccd1 _2426_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3712__A _3712_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3431__B _3437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2328__A _2328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4315__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A2 _3992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2998__A _2998_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__A2 _2420_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__A1 _4268_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__B2 input82/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3515__A1 _4144_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3515__B2 _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2318__A2 _2245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3920__D1 _3331_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2937__S _2937_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output143_A _2125_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3622__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output310_A _2813_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3060__C _3594_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2254__A1 _2254_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2930_ _4320_/Q input56/X _2940_/S vssd1 vssd1 vccd1 vccd1 _3871_/C sky130_fd_sc_hd__mux2_2
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2861_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2888_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2792_ _2799_/A _2812_/B _3378_/C vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__and3_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3219__D _3219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2701__A _2739_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3516__B _4145_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2309__A2 _2424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3413_ _3431_/A _3413_/B _3413_/C vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__or3_1
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2190__B1 _4113_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3344_ _3344_/A vssd1 vssd1 vccd1 vccd1 _4072_/D sky130_fd_sc_hd__clkbuf_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3317_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__A _3564_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2226_ _2226_/A vssd1 vssd1 vccd1 vccd1 _2446_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2478__D1 _2477_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4338__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2493__A1 _2491_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2157_ _2155_/X _2072_/Y _2153_/C _2156_/Y vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__a31oi_2
X_2088_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2529_/A sky130_fd_sc_hd__buf_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1987__A input3/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3993__A1 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2314__C _2414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3745__A1 _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2548__A2 _2547_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3707__A _3707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3426__B _3437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3145__C _3650_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2181__B1 _2180_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3442__A _3457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input139_A spi_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2484__A1 _2287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2236__A1 _2964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3984__A1 _3952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1995__B1 _1942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3736__A1 _2117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3617__A _3617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output260_A _2732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2667__S _2947_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3060_ _3063_/A _3070_/B _3594_/C vssd1 vssd1 vccd1 vccd1 _3061_/A sky130_fd_sc_hd__and3_1
XANTENNA__2894__C _3420_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2011_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2012_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2227__A1 _2225_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3975__A1 _4369_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3962_ _2342_/Y _2357_/A _2357_/Y _3566_/A _3963_/C vssd1 vssd1 vccd1 vccd1 _4363_/D
+ sky130_fd_sc_hd__o2111ai_1
X_2913_ _2913_/A vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2415__B _2557_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1986__B1 _1983_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3893_ _3893_/A _3893_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__and3_1
XANTENNA__4333__D _4333_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2844_ _4305_/Q input40/X _2844_/S vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__mux2_8
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4010__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_9_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3527__A _3564_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2775_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2825_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__2150__B _2182_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4160__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4376_ _4390_/CLK _4376_/D vssd1 vssd1 vccd1 vccd1 _4376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3327_ _3327_/A vssd1 vssd1 vccd1 vccd1 _4066_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2163__B1 _2162_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3262__A _3276_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3258_ _3258_/A vssd1 vssd1 vccd1 vccd1 _4038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2209_ _1968_/Y _3332_/A _1974_/Y _1990_/Y _3301_/A vssd1 vssd1 vccd1 vccd1 _2210_/B
+ sky130_fd_sc_hd__o2111ai_1
X_3189_ _3189_/A vssd1 vssd1 vccd1 vccd1 _4013_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2028__D _2074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3966__A1 _3945_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4243__D _4243_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2044__C _2053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3437__A _3457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2995__B _4230_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2154__B1 _2153_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3172__A _3876_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2457__A1 _2455_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2472__A4 _2445_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2209__A1 _1968_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2235__B _2335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4033__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4153__D _4153_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2950__S _2950_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4183__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3347__A _3347_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput207 _2989_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[9] sky130_fd_sc_hd__buf_2
X_2560_ _2386_/X _2424_/X _4167_/Q vssd1 vssd1 vccd1 vccd1 _2560_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__2251__A _2422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput229 _3143_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput218 _3107_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[18] sky130_fd_sc_hd__buf_2
X_2491_ _4265_/Q vssd1 vssd1 vccd1 vccd1 _2491_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4262_/CLK _4230_/D vssd1 vssd1 vccd1 vccd1 _4230_/Q sky130_fd_sc_hd__dfxtp_1
X_4161_ _4389_/CLK _4161_/D vssd1 vssd1 vccd1 vccd1 _4161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3342__C1 _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3082__A _3082_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2696__A1 input31/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3513__C _3657_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4092_ _4180_/CLK _4092_/D vssd1 vssd1 vccd1 vccd1 _4092_/Q sky130_fd_sc_hd__dfxtp_1
X_3112_ _3239_/C _4205_/Q _3112_/S vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2448__A1 _2448_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3043_ _3186_/B _4186_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3582_/C sky130_fd_sc_hd__mux2_1
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4328__D _4328_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3810__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3945_ _3945_/A _3965_/A _3945_/C _3945_/D vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__and4_1
XANTENNA__2145__B _3294_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2620__A1 _2620_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4063__D _4063_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3876_ _3876_/A vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__buf_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2799__C _3381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2827_ _3215_/B _4092_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _3394_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3257__A _3276_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2758_ _3802_/A _4011_/Q _3790_/A vssd1 vssd1 vccd1 vccd1 _3184_/C sky130_fd_sc_hd__mux2_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2689_ _3893_/A _4049_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _3286_/C sky130_fd_sc_hd__mux2_2
XFILLER_99_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3333__C1 _2155_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4359_ _4390_/CLK _4359_/D vssd1 vssd1 vccd1 vccd1 _4359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2687__A1 input29/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4238__D _4238_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3720__A _3720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4056__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2336__A _2336_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _2061_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2055__B _2055_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2611__A1 _3558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2770__S _3907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3167__A _3192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3317__D _3326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input67_A cpu_sel_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3614__B _3633_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output223_A _3123_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4148__D _4148_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2945__S _2953_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3630__A _3630_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2246__A _2579_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2850__A1 _4026_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3956__B1_N _2306_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _3730_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__nor2_4
XANTENNA__2063__C1 _2059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1991_ _1976_/Y _1977_/X _1986_/Y _1990_/Y vssd1 vssd1 vccd1 vccd1 _2005_/C sky130_fd_sc_hd__o211a_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2602__B2 _2600_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2602__A1 _2281_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3077__A _3081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3661_ _3661_/A _3661_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3662_/A sky130_fd_sc_hd__and3_1
XANTENNA__3158__A2 _2200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2612_ _2581_/X _2582_/X _3996_/A _2579_/X vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__o211a_1
X_3592_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2543_ _2543_/A vssd1 vssd1 vccd1 vccd1 _3369_/A sky130_fd_sc_hd__buf_4
XANTENNA__3563__C1 _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3227__D _3234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3805__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2118__B1 _2117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2474_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__buf_4
X_4213_ _4275_/CLK _4213_/D vssd1 vssd1 vccd1 vccd1 _4213_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2669__A1 input24/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4144_ _4250_/CLK _4144_/D vssd1 vssd1 vccd1 vccd1 _4144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4079__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3243__C _3243_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2855__S _2904_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4058__D _4058_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4075_ _4391_/CLK _4075_/D vssd1 vssd1 vccd1 vccd1 _4075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3026_ _3032_/A _4244_/Q vssd1 vssd1 vccd1 vccd1 _3027_/A sky130_fd_sc_hd__and2_1
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3928_ input16/X _3908_/X _3927_/X _3912_/Y vssd1 vssd1 vccd1 vccd1 _4346_/D sky130_fd_sc_hd__a211o_1
X_3859_ _3859_/A vssd1 vssd1 vccd1 vccd1 _4314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3418__C _3418_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3715__A _3715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3434__B _3459_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3450__A _3450_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input121_A spi_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3085__A1 _4197_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__A1 _4023_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2596__B1 _2595_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2045__C1 _1938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3609__B _3609_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2060__A2 _2152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3328__C _3695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3545__C1 _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3625__A _3625_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2899__A1 _4034_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output173_A _2405_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4221__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3063__C _3596_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2190_ _2129_/A _2129_/B _4113_/Q vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__S _2947_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3360__A _3433_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4371__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3076__A1 _4195_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2704__A _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1974_ _4336_/Q _2659_/A _1971_/Y _1973_/X _1965_/X vssd1 vssd1 vccd1 vccd1 _1974_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3713_ _4242_/Q _3695_/X _3696_/X _3697_/X _3705_/X vssd1 vssd1 vccd1 vccd1 _4242_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3784__C1 _3772_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__B1 _2509_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3644_ _3644_/A _3661_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3645_/A sky130_fd_sc_hd__and3_1
XANTENNA__4341__D _4341_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2339__B1 _2408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3535__A _3546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3575_ _3575_/A vssd1 vssd1 vccd1 vccd1 _4183_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3551__A2 _3536_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2526_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__buf_4
X_2457_ _2455_/Y _2366_/X _2456_/Y vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2388_ _2386_/X _3468_/A _4154_/Q vssd1 vssd1 vccd1 vccd1 _2388_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2511__B1 _2499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2156__A1_N _4068_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4127_ _4177_/CLK _4127_/D vssd1 vssd1 vccd1 vccd1 _4127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3270__A _3270_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4058_ _4326_/CLK _4058_/D vssd1 vssd1 vccd1 vccd1 _4058_/Q sky130_fd_sc_hd__dfxtp_1
X_3009_ _3009_/A vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2290__A2 _2289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2578__B1 _2573_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__C1 _3774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3429__B _3429_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2042__A2 _2018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3148__C _3653_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4251__D _4251_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4244__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3445__A _3953_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3542__A2 _3536_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2502__B1 _2377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3180__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3611__C _3611_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2805__A1 _4088_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2524__A _2579_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output290_A _2879_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2569__B1 _2293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__C1 _3757_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2033__A2 _2141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4161__D _4161_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3518__C1 _3470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__A2 _3764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3355__A _3355_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3533__A2 _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3360_ _3433_/A vssd1 vssd1 vccd1 vccd1 _3381_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3074__B _3089_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2311_ _2517_/A vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__buf_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3291_ _3328_/B _3689_/D _3291_/C _3925_/D vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__and4_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2117_/X _2344_/A _2346_/A _2257_/A _2264_/A vssd1 vssd1 vccd1 vccd1 _2292_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3090__A _3090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2173_ input9/X _2001_/X _2172_/Y _2153_/C vssd1 vssd1 vccd1 vccd1 _2173_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3802__B _3821_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4117__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4336__D _4336_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2434__A _2434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2009__C1 _2137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4267__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2153__B _2153_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1957_ _2022_/A vssd1 vssd1 vccd1 vccd1 _2078_/C sky130_fd_sc_hd__buf_2
XANTENNA__4071__D _4071_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3509__C1 _3504_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2980__B1 _3671_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3627_ _3627_/A vssd1 vssd1 vccd1 vccd1 _4204_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3265__A _3273_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3558_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _4173_/D sky130_fd_sc_hd__nor2_1
X_2509_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__buf_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput118 spi_dat_i[18] vssd1 vssd1 vccd1 vccd1 _2545_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput107 gpio_rty_i vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3489_ _3489_/A vssd1 vssd1 vccd1 vccd1 _3489_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput129 spi_dat_i[28] vssd1 vssd1 vccd1 vccd1 _2620_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3431__C _3431_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4246__D _4246_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2344__A _2344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A3 _2421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__A2 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2971__B1 _3667_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3515__A2 _3308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3175__A _3175_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3920__C1 _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3903__A _3903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3622__B _3635_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2519__A _4267_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4156__D _4156_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2953__S _2953_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output303_A _2939_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2254__A2 _2090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2860_ _2860_/A vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3739__C1 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2791_ _3195_/B _4086_/Q _2937_/S vssd1 vssd1 vccd1 vccd1 _3378_/C sky130_fd_sc_hd__mux2_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2962__A0 _3271_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3516__C _3657_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3412_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3431_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2190__A1 _2129_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3343_ _3343_/A _3343_/B _3343_/C _2069_/Y vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__or4b_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A _3813_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3274_ _3274_/A vssd1 vssd1 vccd1 vccd1 _4045_/D sky130_fd_sc_hd__clkbuf_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2225_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3532__B _3532_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2429__A _2429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2478__C1 _2454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2493__A2 _2411_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _4068_/Q _4070_/Q _3942_/A _2136_/X vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__4066__D _4066_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2087_ _2087_/A vssd1 vssd1 vccd1 vccd1 _2422_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2863__S _2886_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3993__A2 _3992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2989_ _2989_/A vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2314__D _2314_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3745__A2 _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2402__C1 _4390_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2953__A0 _4289_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3426__C _3426_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2181__A1 _4064_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3442__B _3462_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2484__A2 _3468_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2290__B1_N _4148_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2236__A2 _2139_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2641__C1 _2640_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3984__A2 _3955_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1995__A1 _1951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input97_A gpio_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3736__A2 _2539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3109__S _3109_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output253_A _2719_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3633__A _3633_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2172__A1 _1952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2249__A _2382_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3121__A0 _3243_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _4060_/Q _2093_/A _2009_/Y vssd1 vssd1 vccd1 vccd1 _2031_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2227__A2 _2683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _4362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2912_ _2917_/A _2928_/B _3426_/C vssd1 vssd1 vccd1 vccd1 _2913_/A sky130_fd_sc_hd__and3_1
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2415__C _2590_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2632__C1 _2631_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__A2 _3965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1986__A1 _4335_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3892_ _3892_/A vssd1 vssd1 vccd1 vccd1 _4328_/D sky130_fd_sc_hd__clkbuf_1
X_2843_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2872_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2712__A _2712_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2774_ _2774_/A vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3808__A _3808_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3527__B _3527_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2935__A0 _4321_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4305__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4375_ _4390_/CLK _4375_/D vssd1 vssd1 vccd1 vccd1 _4375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2858__S _2858_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3543__A _3546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3326_ _3343_/A _3326_/B _3326_/C _3326_/D vssd1 vssd1 vccd1 vccd1 _3327_/A sky130_fd_sc_hd__or4_1
XANTENNA__2163__A1 _4063_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3262__B _3262_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3112__A0 _3239_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3257_ _3276_/A _3257_/B _3276_/C _3271_/D vssd1 vssd1 vccd1 vccd1 _3258_/A sky130_fd_sc_hd__or4_1
XANTENNA__2159__A _2159_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2208_ _2208_/A vssd1 vssd1 vccd1 vccd1 _2211_/C sky130_fd_sc_hd__inv_2
X_3188_ _3192_/A _3199_/B _3188_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3189_/A sky130_fd_sc_hd__and4_1
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2139_ _2662_/A _3879_/A _2138_/X vssd1 vssd1 vccd1 vccd1 _2139_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3966__A2 _3736_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3718__A _3718_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2622__A _4279_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2044__D _2081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3437__B _3437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2926__A0 _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3453__A _3457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2154__A1 _4071_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2457__A2 _2366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A cpu_adr_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2209__A2 _3332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3628__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4328__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput208 _4394_/A vssd1 vssd1 vccd1 vccd1 gpio_cyc_o sky130_fd_sc_hd__buf_2
Xoutput219 _3111_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[19] sky130_fd_sc_hd__buf_2
X_2490_ _2482_/X _2489_/Y _2404_/X _2469_/X vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__o211a_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4160_ _4172_/CLK _4160_/D vssd1 vssd1 vccd1 vccd1 _4160_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3363__A _3591_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3342__B1 _2153_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3111_ _3111_/A vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__clkbuf_1
X_4091_ _4199_/CLK _4091_/D vssd1 vssd1 vccd1 vccd1 _4091_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2448__A2 _2444_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3042_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3073_/S sky130_fd_sc_hd__buf_2
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2707__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3810__B _3829_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4344__D _4344_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3944_ _2407_/A _2406_/A _3728_/A _2552_/X vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__o22a_1
XANTENNA__2145__C _2145_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3875_ _3875_/A vssd1 vssd1 vccd1 vccd1 _4321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2620__A2 _2628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2826_ _3829_/C _4022_/Q _2826_/S vssd1 vssd1 vccd1 vccd1 _3215_/B sky130_fd_sc_hd__mux2_4
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3257__B _3257_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2757_ _2958_/S vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__buf_4
X_2688_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2954_/S sky130_fd_sc_hd__buf_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3273__A _3273_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__B1 _3805_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4358_ _4390_/CLK _4358_/D vssd1 vssd1 vccd1 vccd1 _4358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A cpu_adr_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3309_ _3309_/A vssd1 vssd1 vccd1 vccd1 _4057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4289_ _4302_/CLK _4289_/D vssd1 vssd1 vccd1 vccd1 _4289_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__D _4254_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A2 _3902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3448__A _3448_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2611__A2 _2526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3167__B _3167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3183__A _3264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3614__C _3624_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_CLK_A clkbuf_2_1_0_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_8_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output216_A _3100_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4150__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__D _4164_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1990_ _4054_/Q _2093_/A _1989_/Y vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2063__B1 _2062_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__A _3470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2602__A2 _2599_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2262__A _3730_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3077__B _3089_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3660_ _3660_/A vssd1 vssd1 vccd1 vccd1 _4218_/D sky130_fd_sc_hd__clkbuf_1
X_2611_ _3558_/B _2526_/A _2606_/Y _2610_/Y vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__o211ai_4
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _3591_/A vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__buf_4
XFILLER_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3563__B1 _3524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2542_ _2406_/X _2407_/X _2408_/X _2409_/X _2541_/Y vssd1 vssd1 vccd1 vccd1 _2542_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3805__B _3805_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3093__A _3099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4212_ _4282_/CLK _4212_/D vssd1 vssd1 vccd1 vccd1 _4212_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2118__A1 _2237_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2473_ _2363_/X _2449_/X _2311_/X _2450_/X _4370_/Q vssd1 vssd1 vccd1 vccd1 _2473_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4143_ _4250_/CLK _4143_/D vssd1 vssd1 vccd1 vccd1 _4143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__D _3260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4339__D _4339_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _4074_/CLK _4074_/D vssd1 vssd1 vccd1 vccd1 _4074_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3821__A _3821_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3025_ _3025_/A vssd1 vssd1 vccd1 vccd1 _3025_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2871__S _2916_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4074__D _4074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2054__B1 _4354_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3268__A _3268_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3927_ _2121_/X _2201_/X _1994_/X _4346_/Q vssd1 vssd1 vccd1 vccd1 _3927_/X sky130_fd_sc_hd__o31a_1
X_3858_ _3871_/A _3877_/B _3858_/C vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__or3_1
X_3789_ _4286_/Q _2200_/A _3748_/A _3736_/Y _3566_/X vssd1 vssd1 vccd1 vccd1 _4286_/D
+ sky130_fd_sc_hd__o221a_1
X_2809_ _3821_/A _4019_/Q _2845_/S vssd1 vssd1 vccd1 vccd1 _3208_/C sky130_fd_sc_hd__mux2_2
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__C _3455_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4023__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4249__D _4249_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3731__A _3765_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4173__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2347__A _3730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input114_A spi_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2045__B1 _2044_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2596__A1 _2526_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3178__A _3192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3609__C _3624_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3328__D _3925_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3545__B1 _2504_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2810__A _3197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output166_A _2318_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4159__D _4159_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__A _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2257__A _2257_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2704__B _4123_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2587__A1 _2526_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1973_ _2055_/B vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__clkbuf_4
X_3712_ _3712_/A vssd1 vssd1 vccd1 vccd1 _4241_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3784__B1 _3771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__B2 _2585_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3643_ _3643_/A vssd1 vssd1 vccd1 vccd1 _4210_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2720__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2339__A1 _2262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3816__A _3816_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3535__B _3535_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3574_ _3574_/A _3584_/B _3657_/A vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__and3_1
XANTENNA__4046__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3551__A3 _3544_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2525_ _2512_/X _2513_/X _3982_/A _2524_/X vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__o211a_1
X_2456_ _2575_/A _2520_/B _2520_/C _2456_/D vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__nand4_2
XFILLER_69_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4069__D _4069_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4126_ _4177_/CLK _4126_/D vssd1 vssd1 vccd1 vccd1 _4126_/Q sky130_fd_sc_hd__dfxtp_1
X_2387_ _2387_/A vssd1 vssd1 vccd1 vccd1 _3468_/A sky130_fd_sc_hd__buf_2
XANTENNA__4196__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2511__A1 _2502_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ _4085_/CLK _4057_/D vssd1 vssd1 vccd1 vccd1 _4057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2167__A _2167_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3008_ _3010_/A _4236_/Q vssd1 vssd1 vccd1 vccd1 _3009_/A sky130_fd_sc_hd__and2_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2578__A1 _3554_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__B1 _2576_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3429__C _3455_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3542__A3 _3528_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2776__S _2825_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3461__A _3461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2502__B2 _2434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2502__A1 _2481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3180__B _3180_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2266__B1 _2117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2569__B2 _2567_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2569__A1 _2281_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__B1 _2541_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4069__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3518__B1 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output283_A _2835_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3636__A _3636_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__A3 _3748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2540__A _2590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3533__A3 _3528_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3074__C _3602_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2310_ _2310_/A1 _2090_/A _2308_/X _2421_/A _2309_/Y vssd1 vssd1 vccd1 vccd1 _3527_/B
+ sky130_fd_sc_hd__a41oi_4
X_3290_ _3707_/A vssd1 vssd1 vccd1 vccd1 _3925_/D sky130_fd_sc_hd__buf_4
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2549__B1_N _4166_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2241_ _4286_/Q _2349_/A _2113_/A vssd1 vssd1 vccd1 vccd1 _2264_/A sky130_fd_sc_hd__o21a_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3371__A _3371_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3802__C _3903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2172_ _1952_/X _2160_/X _4340_/Q vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2715__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2009__B1 _2008_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4352__D _4352_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1956_ _2078_/B vssd1 vssd1 vccd1 vccd1 _1998_/B sky130_fd_sc_hd__buf_2
XANTENNA__2153__C _2153_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3509__B1 _2767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2980__A1 _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3546__A _3546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3626_ _3635_/A _3635_/B _3626_/C vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__or3_1
XANTENNA__2450__A _2450_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3557_ _3557_/A1 _3365_/B _3544_/X _2598_/Y _3547_/X vssd1 vssd1 vccd1 vccd1 _4172_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3265__B _3279_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2508_ _2506_/Y _2411_/X _2507_/Y vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__o21a_4
Xinput108 spi_ack_i vssd1 vssd1 vccd1 vccd1 _2384_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3488_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput119 spi_dat_i[19] vssd1 vssd1 vccd1 vccd1 _3551_/A1 sky130_fd_sc_hd__buf_2
X_2439_ _4260_/Q vssd1 vssd1 vccd1 vccd1 _2439_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3281__A _3297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2496__B1 _2495_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4109_ _4251_/CLK _4109_/D vssd1 vssd1 vccd1 vccd1 _4109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4211__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4262__D _4262_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3456__A _3456_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2971__A1 _2197_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4361__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_25_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3920__B1 _2008_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input42_A cpu_dat_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3191__A _3191_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3684__C1 _3683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3622__C _3622_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2239__B1 _2238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2254__A3 _2248_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3987__B1 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4172__D _4172_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3739__B1 _3735_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2790_ _3815_/C _4016_/Q _2826_/S vssd1 vssd1 vccd1 vccd1 _3195_/B sky130_fd_sc_hd__mux2_2
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3366__A _3366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2962__A1 _4218_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_16_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4282_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2270__A _2367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3411_ _3411_/A vssd1 vssd1 vccd1 vccd1 _4099_/D sky130_fd_sc_hd__clkbuf_1
X_4391_ _4391_/CLK _4391_/D vssd1 vssd1 vccd1 vccd1 _4391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3342_ _4071_/Q _3314_/A _2153_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _4071_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3911__B1 _4336_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2190__A2 _2129_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B _3821_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3273_ _3273_/A _3279_/B _3273_/C _3286_/D vssd1 vssd1 vccd1 vccd1 _3274_/A sky130_fd_sc_hd__and4_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2478__B1 _2453_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2224_ _2328_/A vssd1 vssd1 vccd1 vccd1 _2224_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2155_ _1971_/C _1971_/D _1998_/B _4348_/Q vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4347__D _4347_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4234__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2086_ _2129_/A _2106_/A _4146_/Q vssd1 vssd1 vccd1 vccd1 _2087_/A sky130_fd_sc_hd__o21bai_2
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2445__A _2531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1989__C1 _1977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4082__D _4082_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4384__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2988_ _2988_/A _4227_/Q vssd1 vssd1 vccd1 vccd1 _2989_/A sky130_fd_sc_hd__and2_1
XANTENNA__3745__A3 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2402__B1 _2429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3276__A _3276_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1939_ input8/X vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2953__A1 input69/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput90 gpio_dat_i[24] vssd1 vssd1 vccd1 vccd1 _2590_/D sky130_fd_sc_hd__clkbuf_2
X_3609_ _3609_/A _3609_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3610_/A sky130_fd_sc_hd__and3_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2181__A2 _1977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3442__C _3442_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4257__D _4257_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2641__B1 _2636_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2074__B _2081_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1995__A2 _1994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3186__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2090__A _2090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4107__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3914__A _3914_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output246_A _2217_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3633__B _3633_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2172__A2 _2160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2249__B _2383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4167__D _4167_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4257__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3121__A1 _4207_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4390_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2880__A0 _4311_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2265__A _2453_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3960_ _3960_/A _3973_/B _3963_/C vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__and3_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2911_ _3250_/B _4106_/Q _2911_/S vssd1 vssd1 vccd1 vccd1 _3426_/C sky130_fd_sc_hd__mux2_1
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2415__D _2415_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2632__B1 _2509_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1986__A2 _2182_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3891_ _3895_/A _3935_/B _3891_/C vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__or3_1
X_2842_ _2842_/A vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2773_ _2799_/A _2780_/B _3372_/A vssd1 vssd1 vccd1 vccd1 _2774_/A sky130_fd_sc_hd__and3_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3096__A _3099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2935__A1 input58/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3824__A _3824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2699__B1 _3466_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4374_ _4380_/CLK _4374_/D vssd1 vssd1 vccd1 vccd1 _4374_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3543__B _3543_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3325_ _4065_/Q _3314_/A _2184_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _4065_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2163__A2 _2093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3262__C _3276_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3256_ _3295_/C vssd1 vssd1 vccd1 vccd1 _3276_/C sky130_fd_sc_hd__clkbuf_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__D _4077_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3112__A1 _4205_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2159__B _2159_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2207_ _2207_/A _2207_/B _2207_/C _2207_/D vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__nand4_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3187_ _3187_/A vssd1 vssd1 vccd1 vccd1 _4012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2871__A0 _3234_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2138_ _2136_/X _3942_/A _4043_/Q vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1998__B _1998_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2069_ _2134_/A _3935_/C _2068_/X vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2175__A _2175_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3966__A3 _2255_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2903__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3437__C _3437_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2926__A1 _4039_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3734__A _3767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3453__B _3462_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2154__A2 _2093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2784__S _3907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2862__A0 _4308_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2085__A _2085_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2614__B1 _2613_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3909__A _3945_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2813__A _2813_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output196_A _3031_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput209 _3041_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__2959__S _3161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3644__A _3644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3342__A1 _4071_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3110_ _3117_/A _3125_/B _3626_/C vssd1 vssd1 vccd1 vccd1 _3111_/A sky130_fd_sc_hd__and3_1
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ _4251_/CLK _4090_/D vssd1 vssd1 vccd1 vccd1 _4090_/Q sky130_fd_sc_hd__dfxtp_1
X_3041_ _3041_/A vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2694__S _3161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2448__A3 _2308_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3810__C _3810_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2707__B _4124_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2605__B1 _2604_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _4356_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2145__D _2145_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2723__A _2723_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3874_ _3874_/A _3893_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__and3_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3819__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2620__A3 _2514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2825_ _4302_/Q input37/X _2825_/S vssd1 vssd1 vccd1 vccd1 _3829_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4360__D _4360_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3257__C _3276_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2756_ _4291_/Q input35/X _3907_/A vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3554__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2869__S _2905_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2687_ _4329_/Q input29/X _2953_/S vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3273__B _3279_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__A1 _2201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4357_ _4391_/CLK _4357_/D vssd1 vssd1 vccd1 vccd1 _4357_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3308_/A _3774_/A _3308_/C vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__and3_1
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4326_/CLK _4288_/D vssd1 vssd1 vccd1 vccd1 _4288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3239_ _3247_/A _3253_/B _3239_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3240_/A sky130_fd_sc_hd__and4_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2844__A0 _4305_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3729__A _3764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4270__D _4270_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3167__C _3167_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2779__S _2937_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3464__A _3800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3088__A0 _3219_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output209_A _3041_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2543__A _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3639__A _3639_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2063__A1 _2061_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3358__B _3365_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4180__D _4180_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3077__C _3605_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2610_ _2474_/X _2452_/X _2453_/X _2454_/X _2609_/Y vssd1 vssd1 vccd1 vccd1 _2610_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3590_ _3590_/A vssd1 vssd1 vccd1 vccd1 _4189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3563__A1 _4178_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3563__B2 _2644_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2541_ _2538_/Y _3617_/A _2540_/Y vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__2689__S _2954_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3374__A _3383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2472_ _2472_/A1 _2444_/X _2308_/X _2445_/X _2471_/Y vssd1 vssd1 vccd1 vccd1 _3541_/B
+ sky130_fd_sc_hd__a41oi_4
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3805__C _3805_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3093__B _3106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2118__A2 _2393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4211_ _4275_/CLK _4211_/D vssd1 vssd1 vccd1 vccd1 _4211_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2523__C1 _2522_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ _4250_/CLK _4142_/D vssd1 vssd1 vccd1 vccd1 _4142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2718__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4073_ _4085_/CLK _4073_/D vssd1 vssd1 vccd1 vccd1 _4073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3821__B _3821_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3024_ _3032_/A _4243_/Q vssd1 vssd1 vccd1 vccd1 _3025_/A sky130_fd_sc_hd__and2_1
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2826__A0 _3829_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4355__D _4355_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3549__A _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2453__A _2453_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2054__A1 _1952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3926_ _3926_/A vssd1 vssd1 vccd1 vccd1 _4345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4090__D _4090_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3857_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3877_/B sky130_fd_sc_hd__clkbuf_2
X_3788_ _4285_/Q _2133_/A _2407_/X _2406_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4285_/D
+ sky130_fd_sc_hd__o221a_1
X_2808_ _4299_/Q input65/X _2844_/S vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__mux2_8
X_2739_ _2739_/A vssd1 vssd1 vccd1 vccd1 _2748_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3284__A _3284_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2628__A _2628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2817__A0 _3210_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4318__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4265__D _4265_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A gpio_rty_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2363__A _2452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3459__A _3459_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2045__A1 _4344_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2596__A2 _3556_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3178__B _3199_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3545__A1 _2503_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input72_A cpu_we_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3194__A _3343_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output159_A _2588_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2538__A _4269_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2808__A0 _4299_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4175__D _4175_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3369__A _3369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2273__A _2336_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ _1951_/A _1994_/A _2201_/A vssd1 vssd1 vccd1 vccd1 _2055_/B sky130_fd_sc_hd__o21bai_4
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3711_ _3717_/A _4241_/Q _3721_/C _3711_/D vssd1 vssd1 vccd1 vccd1 _3712_/A sky130_fd_sc_hd__and4_1
XANTENNA__3784__A1 _4282_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3784__B2 input98/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__A2 _2584_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3642_ _3659_/A _3659_/B _3642_/C vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__or3_1
XANTENNA__2339__A2 _2375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2720__B _4130_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3573_ _3573_/A vssd1 vssd1 vccd1 vccd1 _4182_/D sky130_fd_sc_hd__clkbuf_1
X_2524_ _2579_/A vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2455_ _4261_/Q vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2386_ _2644_/A vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__buf_2
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3832__A _3832_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4125_ _4177_/CLK _4125_/D vssd1 vssd1 vccd1 vccd1 _4125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2511__A2 _2510_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3043__S _3073_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _4074_/CLK _4056_/D vssd1 vssd1 vccd1 vccd1 _4056_/Q sky130_fd_sc_hd__dfxtp_1
X_3007_ _3007_/A vssd1 vssd1 vccd1 vccd1 _3007_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3472__B1 _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2882__S _2916_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4085__D _4085_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3279__A _3328_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3775__A1 _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2578__A2 _2362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3909_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3909_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_7_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4140__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2502__A2 _2501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3180__C _3195_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4290__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2266__A1 _2367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3189__A _3189_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2093__A _2093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2569__A2 _2566_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__A1 _3752_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3518__A1 _2225_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output276_A _2699_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2540__B _2557_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3128__S _3147_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__D1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2099_/Y _2964_/A _2393_/A vssd1 vssd1 vccd1 vccd1 _2344_/A sky130_fd_sc_hd__a21boi_4
XANTENNA__3652__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2268__A _4251_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2171_ _4060_/Q vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2715__B _4128_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3099__A _3099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2009__A1 _2006_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1955_ _4357_/Q _2201_/A vssd1 vssd1 vccd1 vccd1 _2078_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4013__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2731__A _2737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3827__A _3827_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3509__B2 _3490_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3509__A1 _4140_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3546__B _3546_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2980__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4163__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3625_ _3625_/A vssd1 vssd1 vccd1 vccd1 _4203_/D sky130_fd_sc_hd__clkbuf_1
X_3556_ _3558_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _4171_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3265__C _3265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2507_ _2507_/A _2557_/B _2507_/C _2507_/D vssd1 vssd1 vccd1 vccd1 _2507_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__2877__S _2911_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput109 spi_dat_i[0] vssd1 vssd1 vccd1 vccd1 _2254_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_3487_ _3487_/A vssd1 vssd1 vccd1 vccd1 _4129_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3562__A _3562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2438_ _3536_/A _2436_/X _2437_/Y vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_97_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2496__A1 _2496_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2369_ _2365_/Y _2366_/X _2368_/Y vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4284_/CLK _4108_/D vssd1 vssd1 vccd1 vccd1 _4108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4039_ _4225_/CLK _4039_/D vssd1 vssd1 vccd1 vccd1 _4039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2462__A_N _2382_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2971__A2 _2200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3920__A1 _2006_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3684__B1 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2088__A _2422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input35_A cpu_dat_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2239__A1 _3578_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3987__B2 _2563_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3987__A1 _3968_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4036__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2254__A4 _2421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3739__A1 _4252_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3739__B2 input85/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3647__A _3647_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4186__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3410_ _3410_/A _3429_/B _3424_/C vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__and3_1
X_4390_ _4390_/CLK _4390_/D vssd1 vssd1 vccd1 vccd1 _4390_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2697__S _2954_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3341_ _4070_/Q _3331_/X _3340_/X _3346_/C vssd1 vssd1 vccd1 vccd1 _4070_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3911__A1 _2121_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3382__A _3382_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3272_ _3272_/A vssd1 vssd1 vccd1 vccd1 _4044_/D sky130_fd_sc_hd__clkbuf_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__C _3831_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2223_ _2581_/A vssd1 vssd1 vccd1 vccd1 _2328_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2478__A1 _2474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2154_ _4071_/Q _2093_/X _2153_/Y vssd1 vssd1 vccd1 vccd1 _2158_/B sky130_fd_sc_hd__o21ai_1
XFILLER_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2726__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2085_ _2085_/A _2085_/B _2085_/C _2085_/D vssd1 vssd1 vccd1 vccd1 _2106_/A sky130_fd_sc_hd__nand4_4
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4363__D _4363_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1989__B1 _1988_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2987_ _2987_/A vssd1 vssd1 vccd1 vccd1 _2987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2402__B2 _2434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2402__A1 _3730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1938_ _1938_/A vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__buf_2
XANTENNA__3276__B _3276_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput91 gpio_dat_i[25] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_2
Xinput80 gpio_dat_i[15] vssd1 vssd1 vccd1 vccd1 _2507_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ _3608_/A vssd1 vssd1 vccd1 vccd1 _4196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2166__B1 _2165_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ _3546_/A _3539_/B vssd1 vssd1 vccd1 vccd1 _4157_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3292__A _3292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4059__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2641__A1 _3562_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4273__D _4273_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2074__C _2081_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3467__A _3467_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3186__B _3186_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2157__B1 _2156_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3914__B _3942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3633__C _3648_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output239_A _3071_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3141__S _3147_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2880__A1 input47/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2632__A1 _2526_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4183__D _4183_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2910_ _3863_/C _4036_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _3250_/B sky130_fd_sc_hd__mux2_4
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2632__B2 _2630_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3890_ _3890_/A vssd1 vssd1 vccd1 vccd1 _4327_/D sky130_fd_sc_hd__clkbuf_1
X_2841_ _2859_/A _2841_/B _3398_/C vssd1 vssd1 vccd1 vccd1 _2842_/A sky130_fd_sc_hd__and3_1
XANTENNA__3377__A _3377_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2281__A _2380_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2772_ _3188_/C _4083_/Q _2955_/S vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3096__B _3106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3345__C1 _3315_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2148__B1 _2078_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2699__A1 _2677_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4373_ _4391_/CLK _4373_/D vssd1 vssd1 vccd1 vccd1 _4373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3324_ _3324_/A vssd1 vssd1 vccd1 vccd1 _4064_/D sky130_fd_sc_hd__clkbuf_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4358__D _4358_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4201__CLK _4201_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3262__D _3271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3255_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3840__A _3840_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2206_ _2662_/A _3914_/A _2205_/Y vssd1 vssd1 vccd1 vccd1 _2207_/C sky130_fd_sc_hd__o21ai_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3195_/A _3186_/B _3195_/C _3190_/D vssd1 vssd1 vccd1 vccd1 _3187_/A sky130_fd_sc_hd__or4_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3051__S _3073_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2456__A _2575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2871__A1 _4099_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2137_ _2137_/A vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1998__C _2053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4351__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _2055_/A _2055_/B _4072_/Q vssd1 vssd1 vccd1 vccd1 _2068_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2175__B _2175_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4093__D _4093_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3966__A4 _3724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3287__A _3287_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2139__B1 _2138_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3453__C _3453_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4268__D _4268_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3750__A _3767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input137_A spi_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2366__A _2366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2862__A1 input43/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2085__B _2085_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2075__C1 _1938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2614__A1 _3559_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3197__A _3197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output189_A _3016_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__A _3940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4224__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3644__B _3661_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2425__B1_N _4155_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3342__A2 _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2975__S _3150_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2550__B1 _2549_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__D _4178_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3660__A _3660_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4374__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3040_ _3044_/A _3052_/B _3580_/A vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__and3_1
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2448__A4 _2445_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2605__A1 _2605_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3942_ _3942_/A _3942_/B _3942_/C vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__and3_1
X_3873_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3819__B _3829_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2824_ _2824_/A vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2620__A4 _2531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2369__B1 _2368_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3257__D _3271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3835__A _3835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2755_ _2957_/S vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__clkbuf_4
X_2686_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2953_/S sky130_fd_sc_hd__buf_4
XANTENNA__3554__B _3554_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4356_ _4356_/CLK _4356_/D vssd1 vssd1 vccd1 vccd1 _4356_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3273__C _3273_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__A2 input18/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4088__D _4088_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2541__B1 _2540_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3307_ _3433_/A vssd1 vssd1 vccd1 vccd1 _3774_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2885__S _2885_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3570__A _3570_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4287_ _4302_/CLK _4287_/D vssd1 vssd1 vccd1 vccd1 _4287_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3238_ _3264_/A vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ input1/X vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__inv_2
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2844__A1 input40/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4247__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3557__C1 _3547_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3167__D _3945_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2532__B1 _2530_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2795__S _2844_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3480__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3088__A1 _4198_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2824__A _2824_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2599__B1 _2598_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2063__A2 _2001_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__C _3358_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3548__C1 _3547_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3655__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2540_ _2590_/A _2557_/B _2590_/C _2540_/D vssd1 vssd1 vccd1 vccd1 _2540_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__3563__A2 _3447_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3374__B _3389_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2471_ _2330_/X _2446_/X _4159_/Q vssd1 vssd1 vccd1 vccd1 _2471_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2771__A0 _3807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3093__C _3614_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4210_ _4282_/CLK _4210_/D vssd1 vssd1 vccd1 vccd1 _4210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2523__B1 _2518_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4141_ _4141_/CLK _4141_/D vssd1 vssd1 vccd1 vccd1 _4141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3390__A _3390_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2718__B _4129_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4072_ _4085_/CLK _4072_/D vssd1 vssd1 vccd1 vccd1 _4072_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3821__C _3831_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3023_ _3023_/A vssd1 vssd1 vccd1 vccd1 _3032_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2826__A1 _4022_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2734__A _2734_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3787__C1 _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2054__A2 _2160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3925_ _3940_/C _3925_/B _3925_/C _3925_/D vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__and4_1
XANTENNA__4371__D _4371_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3856_ _3856_/A vssd1 vssd1 vccd1 vccd1 _4313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2807_ _2807_/A vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__clkbuf_1
X_3787_ _2117_/X _3586_/B _3729_/X _3732_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4284_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3565__A _3724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2738_ _2738_/A vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2669_ _4326_/Q input24/X _2949_/S vssd1 vssd1 vccd1 vccd1 _3887_/C sky130_fd_sc_hd__mux2_2
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4339_ _4347_/CLK _4339_/D vssd1 vssd1 vccd1 vccd1 _4339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2628__B _2644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2278__C1 _2277_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2817__A1 _4090_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2644__A _2644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3459__B _3459_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2045__A2 _1970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4281__D _4281_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3178__C _3178_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3475__A _3475_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3545__A2 _3536_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input65_A cpu_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2505__B1 _2504_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2819__A _2819_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output221_A _3114_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2808__A1 input65/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3710_ _4240_/Q _3695_/X _3696_/X _3697_/X _3705_/X vssd1 vssd1 vccd1 vccd1 _4240_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4191__D _4191_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1971_ input5/X _1998_/B _1971_/C _1971_/D vssd1 vssd1 vccd1 vccd1 _1971_/Y sky130_fd_sc_hd__nand4b_2
XANTENNA__3784__A2 _3657_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3659_/B sky130_fd_sc_hd__clkbuf_2
X_3572_ _3586_/A _3586_/B _3572_/C vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__or3_1
XANTENNA__3385__A _3433_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2523_ _3546_/B _2362_/X _2518_/Y _2522_/Y vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__o211ai_4
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2454_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2385_ _2382_/X _2383_/X _2385_/C _2503_/D vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__2729__A _2737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4124_ _4177_/CLK _4124_/D vssd1 vssd1 vccd1 vccd1 _4124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4366__D _4366_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 RST_N vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _4302_/CLK _4055_/D vssd1 vssd1 vccd1 vccd1 _4055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3006_ _3010_/A _4235_/Q vssd1 vssd1 vccd1 vccd1 _3007_/A sky130_fd_sc_hd__and2_1
XANTENNA__3472__A1 _2739_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3279__B _3279_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3775__A2 _3764_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2983__A0 _3291_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__clkbuf_2
X_3839_ _3847_/A _3853_/B _3839_/C vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__or3_1
XANTENNA__3295__A _3591_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3160__B1 _3576_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4276__D _4276_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3180__D _3190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2266__A2 _2335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3766__A2 _3764_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3518__A2 _3308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2540__C _2590_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output269_A _2672_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__C1 _3909_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output171_A _2359_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3144__S _3144_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4186__D _4186_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2170_ _4062_/Q _1977_/X _2169_/Y vssd1 vssd1 vccd1 vccd1 _2175_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__2983__S _3157_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2284__A _2284_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3099__B _3106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2009__A2 _2168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1954_ input6/X vssd1 vssd1 vccd1 vccd1 _1961_/A sky130_fd_sc_hd__clkinv_2
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2731__B _4135_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3509__A2 _3308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3624_ _3624_/A _3633_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__and3_1
XANTENNA__4308__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ _4170_/Q _3447_/A _3524_/X _2583_/X _3547_/X vssd1 vssd1 vccd1 vccd1 _4170_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3843__A _3847_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3265__D _3286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3486_ _3492_/A _4129_/Q _3502_/C vssd1 vssd1 vccd1 vccd1 _3487_/A sky130_fd_sc_hd__and3_1
X_2506_ _4266_/Q vssd1 vssd1 vccd1 vccd1 _2506_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2437_ _2287_/X _3468_/A _4156_/Q vssd1 vssd1 vccd1 vccd1 _2437_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__3562__B _3562_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2496__A2 _2420_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2368_ _2575_/A _2520_/B _2520_/C _2368_/D vssd1 vssd1 vccd1 vccd1 _2368_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__2350__D1 _3744_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4096__D _4096_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2299_ _4252_/Q _2295_/X _2298_/X input85/X vssd1 vssd1 vccd1 vccd1 _2299_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2893__S _2916_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4107_ _4286_/CLK _4107_/D vssd1 vssd1 vccd1 vccd1 _4107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4038_ _4085_/CLK _4038_/D vssd1 vssd1 vccd1 vccd1 _4038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2405__C1 _2373_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2956__B1 _3361_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3920__A2 _3902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput190 _3018_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3684__B2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__A1 _4228_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A cpu_adr_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2239__A2 _2236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3987__A2 _3969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3739__A2 _3734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2947__A0 _3167_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1972__B1_N _2201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3340_ _4350_/Q _3907_/A _2074_/Y _3805_/B vssd1 vssd1 vccd1 vccd1 _3340_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3911__A2 _2201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3663__A _3804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3124__A0 _3245_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3271_ _3276_/A _3271_/B _3276_/C _3271_/D vssd1 vssd1 vccd1 vccd1 _3272_/A sky130_fd_sc_hd__or4_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2452_/A _3730_/B _2429_/A _2552_/A _4390_/Q vssd1 vssd1 vccd1 vccd1 _2581_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__2478__A2 _2452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _2153_/A _2153_/B _2153_/C vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__nand3_1
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2726__B _4133_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_6_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2084_ _2084_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2085_/D sky130_fd_sc_hd__nor2_1
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1989__A1 _1987_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2742__A _2748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4130__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3838__A _3838_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2986_ _2988_/A _4226_/Q vssd1 vssd1 vccd1 vccd1 _2987_/A sky130_fd_sc_hd__and2_1
XANTENNA__2402__A2 _2428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1937_ _4058_/Q _2184_/C _1936_/Y vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__3276__C _3276_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput81 gpio_dat_i[16] vssd1 vssd1 vccd1 vccd1 _2520_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4280__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3607_ _3611_/A _3611_/B _3607_/C vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__or3_1
Xinput70 cpu_sel_i[3] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_4
Xinput92 gpio_dat_i[26] vssd1 vssd1 vccd1 vccd1 _2608_/D sky130_fd_sc_hd__clkbuf_2
X_3538_ _2436_/C _3536_/X _3528_/X _2437_/Y _3537_/X vssd1 vssd1 vccd1 vccd1 _4156_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3573__A _3573_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2166__A1 _4061_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3469_ _3490_/A vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__buf_2
XANTENNA__2189__A _2683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2917__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2626__C1 _2625_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2641__A2 _2526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3748__A _3748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2074__D _2074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3186__C _3195_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2798__S _2955_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3483__A _3935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2157__A1 _2155_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3914__C _3914_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2099__A _4250_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output301_A _2934_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2617__C1 _2616_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4153__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3658__A _3658_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2840_ _3219_/B _4094_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _3398_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2632__A2 _2629_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2771_ _3807_/A _4013_/Q _3790_/A vssd1 vssd1 vccd1 vccd1 _3188_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3096__C _3618_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3393__A _3441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3345__B1 _2059_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2148__A1 _4349_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2699__A2 _2680_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4372_ _4390_/CLK _4372_/D vssd1 vssd1 vccd1 vccd1 _4372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3323_ _3343_/A _3326_/C _3323_/C _2186_/C vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__or4b_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3254_/A vssd1 vssd1 vccd1 vccd1 _4037_/D sky130_fd_sc_hd__clkbuf_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _3942_/C _1996_/X _1949_/Y vssd1 vssd1 vccd1 vccd1 _2205_/Y sky130_fd_sc_hd__o21ai_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2737__A _2737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2320__A1 _2319_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3185_ _3185_/A vssd1 vssd1 vccd1 vccd1 _4011_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2456__B _2520_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1998__D _2081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2136_ _2136_/A vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__buf_2
XANTENNA__4374__D _4374_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2067_ _2065_/Y _2001_/A _2066_/Y vssd1 vssd1 vccd1 vccd1 _3935_/C sky130_fd_sc_hd__o21ai_2
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2175__C _2175_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3568__A _3720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _2197_/X _2200_/X _3664_/C vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2139__A1 _2662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4026__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4176__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4284__D _4284_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2075__B1 _2074_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2085__C _2085_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2382__A _2382_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3478__A _3478_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2614__A2 _2420_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input95_A gpio_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3925__B _3925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3644__C _3648_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output251_A _2714_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2550__A1 _3551_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3941__A _3941_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2557__A _2590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4194__D _4194_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2066__B1 _4352_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2605__A2 _2444_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3388__A _3461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3941_ _3941_/A vssd1 vssd1 vccd1 vccd1 _4355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2292__A _2292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3872_ _3872_/A vssd1 vssd1 vccd1 vccd1 _4320_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3819__C _3819_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2823_ _2828_/A _2841_/B _3391_/A vssd1 vssd1 vccd1 vccd1 _2824_/A sky130_fd_sc_hd__and3_1
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2754_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2369__A1 _2365_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4049__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2685_ _2677_/X _2680_/X _3457_/C vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__o21a_2
XFILLER_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4369__D _4369_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4199__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4355_ _4391_/CLK _4355_/D vssd1 vssd1 vccd1 vccd1 _4355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3273__D _3286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__A3 _1918_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2541__A1 _2538_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3306_ _3953_/C vssd1 vssd1 vccd1 vccd1 _3433_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3851__A _3851_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4286_ _4286_/CLK _4286_/D vssd1 vssd1 vccd1 vccd1 _4286_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3062__S _3076_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3237_ _3237_/A vssd1 vssd1 vccd1 vccd1 _4030_/D sky130_fd_sc_hd__clkbuf_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ _3168_/A vssd1 vssd1 vccd1 vccd1 _4007_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2186__B _2186_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2119_ _2346_/A _2257_/A _2517_/A _2450_/A vssd1 vssd1 vccd1 vccd1 _2357_/A sky130_fd_sc_hd__o22ai_4
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3099_ _3099_/A _3106_/B _3620_/A vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__and3_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3298__A _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3557__B1 _2598_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4279__D _4279_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2532__A1 _3466_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2532__B2 _3544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__B _4127_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2377__A _3728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A cpu_adr_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2599__A1 _3557_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3001__A _3023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output299_A _2924_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3548__B1 _3524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3936__A _3936_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3655__B _3659_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3147__S _3147_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3374__C _3374_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2470_ _2461_/X _2468_/Y _2404_/X _2469_/X vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2771__A1 _4013_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4341__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4189__D _4189_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4140_ _4141_/CLK _4140_/D vssd1 vssd1 vccd1 vccd1 _4140_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2523__A1 _3546_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3671__A _3671_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2287__A _2529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _4074_/CLK _4071_/D vssd1 vssd1 vccd1 vccd1 _4071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3022_ _3022_/A vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3484__C1 _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3787__B1 _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3924_ _2044_/A _3902_/X _2179_/Y _3566_/A _3331_/X vssd1 vssd1 vccd1 vccd1 _4344_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2750__A _2752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3846__A _3846_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3855_ _3855_/A _3869_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__and3_1
X_2806_ _2828_/A _2812_/B _3383_/C vssd1 vssd1 vccd1 vccd1 _2807_/A sky130_fd_sc_hd__and3_2
X_3786_ _3734_/X _2236_/X _2238_/X _3938_/D _2398_/X vssd1 vssd1 vccd1 vccd1 _4283_/D
+ sky130_fd_sc_hd__o2111a_1
X_2737_ _2737_/A _4138_/Q vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__and2_1
XANTENNA__2471__B1_N _4159_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2668_ _2128_/X _2133_/X _3451_/A vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4099__D _4099_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2599_ _3557_/A1 _2420_/X _2421_/X _2598_/Y vssd1 vssd1 vccd1 vccd1 _2599_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__3581__A _3581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4338_ _4347_/CLK _4338_/D vssd1 vssd1 vccd1 vccd1 _4338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2197__A _3036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _4280_/CLK _4269_/D vssd1 vssd1 vccd1 vccd1 _4269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A cpu_adr_i[0] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2628__C _2628_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2278__B1 _2261_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4214__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2644__B _2644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__B1 _3771_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3459__C _3466_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3178__D _3945_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4364__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2660__A _2957_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3545__A3 _3544_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2202__B1 _4337_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input58_A cpu_dat_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2505__A1 _2283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2835__A _2835_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output214_A _3094_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ _1970_/A vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2441__B1 _2440_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3666__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3640_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__clkbuf_2
X_3571_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__clkbuf_2
X_2522_ _2474_/X _2452_/X _2453_/X _2454_/X _2521_/Y vssd1 vssd1 vccd1 vccd1 _2522_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2453_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2729__B _4134_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2384_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _4172_/CLK _4123_/D vssd1 vssd1 vccd1 vccd1 _4123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 cpu_adr_i[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
X_4054_ _4326_/CLK _4054_/D vssd1 vssd1 vccd1 vccd1 _4054_/Q sky130_fd_sc_hd__dfxtp_1
X_3005_ _3005_/A vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4237__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2745__A _2745_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3472__A2 _2248_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4387__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4382__D _4382_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3279__C _3279_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3576__A _3586_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__B1 _2431_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__A3 _3765_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2983__A1 _4225_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3838_ _3838_/A vssd1 vssd1 vccd1 vccd1 _4305_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3295__B _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3932__B1 _4350_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3160__A1 _2988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input112_A spi_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2671__A0 _3276_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__D _4292_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3486__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__A3 _3765_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2390__A _4258_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4347_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2540__D _2540_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__B1 _2024_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output164_A _2627_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3099__C _3620_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3396__A _3396_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1953_ _1952_/X _1932_/X _4337_/Q vssd1 vssd1 vccd1 vccd1 _1962_/B sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_19_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4286_/CLK sky130_fd_sc_hd__clkbuf_16
X_3623_ _3623_/A vssd1 vssd1 vccd1 vccd1 _4202_/D sky130_fd_sc_hd__clkbuf_1
X_3554_ _3558_/A _3554_/B vssd1 vssd1 vccd1 vccd1 _4169_/D sky130_fd_sc_hd__nor2_1
X_3485_ _3976_/A vssd1 vssd1 vccd1 vccd1 _3502_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_2505_ _2283_/X _2503_/X _2504_/Y vssd1 vssd1 vccd1 vccd1 _2505_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3843__B _3853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2436_ _2382_/X _2383_/X _2436_/C _2503_/D vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4377__D _4377_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2496__A3 _2421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2350__C1 _2414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2367_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2575_/A sky130_fd_sc_hd__buf_2
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2298_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2298_/X sky130_fd_sc_hd__buf_4
X_4106_ _4180_/CLK _4106_/D vssd1 vssd1 vccd1 vccd1 _4106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2475__A _4263_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4037_ _4199_/CLK _4037_/D vssd1 vssd1 vccd1 vccd1 _4037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2405__B1 _2404_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2956__A1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2169__C1 _2153_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput180 _2998_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput191 _3020_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__4287__D _4287_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__A2 _3351_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2341__C1 _2125_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2892__A0 _3855_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2947__A1 _4077_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output281_A _2824_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2240__B1_N _2393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4082__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3911__A3 _1994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3155__S _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2580__C1 _2579_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3270_ _3270_/A vssd1 vssd1 vccd1 vccd1 _4043_/D sky130_fd_sc_hd__clkbuf_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3124__A1 _4208_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2221_ _2450_/A vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4197__D _4197_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2152_ _2152_/A vssd1 vssd1 vccd1 vccd1 _2153_/C sky130_fd_sc_hd__buf_2
XANTENNA__2295__A _3720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2083_ _2083_/A _2083_/B _2083_/C _2083_/D vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__nand4_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2635__B1 _2634_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1989__A2 _2168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2742__B _4140_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2985_ _3023_/A vssd1 vssd1 vccd1 vccd1 _2988_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1936_ _3916_/B _3916_/C _1977_/A vssd1 vssd1 vccd1 vccd1 _1936_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3854__A _3854_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3276__D _3317_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput82 gpio_dat_i[17] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_2
X_3606_ _3606_/A vssd1 vssd1 vccd1 vccd1 _4195_/D sky130_fd_sc_hd__clkbuf_1
Xinput71 cpu_stb_i vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__clkbuf_4
Xinput60 cpu_dat_i[3] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_4
Xinput93 gpio_dat_i[27] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
X_3537_ _3547_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2166__A2 _1977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3468_ _3468_/A vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2419_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__clkbuf_2
X_3399_ _3399_/A vssd1 vssd1 vccd1 vccd1 _4094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2917__B _2928_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2626__B1 _2621_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2933__A _2943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3051__A0 _3190_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3764__A _3764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3186__D _3190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2157__A2 _2072_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2562__C1 _4378_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input40_A cpu_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2865__A0 _3231_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3004__A _3010_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2617__B1 _2509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2843__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2770_ _4293_/Q input57/X _3907_/A vssd1 vssd1 vccd1 vccd1 _3807_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3674__A _3674_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3345__A1 _4073_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2148__A2 _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2553__C1 _4377_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4371_ _4371_/CLK _4371_/D vssd1 vssd1 vccd1 vccd1 _4371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3322_ _4063_/Q _3314_/X _2162_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _4063_/D sky130_fd_sc_hd__o211a_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3273_/A _3253_/B _3253_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3254_/A sky130_fd_sc_hd__and4_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2305__C1 _4359_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2204_ _2204_/A vssd1 vssd1 vccd1 vccd1 _3942_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__1922__A _4356_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3184_ _3192_/A _3199_/B _3184_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3185_/A sky130_fd_sc_hd__and4_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2737__B _4138_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2320__A2 _2289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2135_ _4323_/Q input72/X _2659_/A vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_4
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2456__C _2520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2066_ _1952_/A _2160_/A _4352_/Q vssd1 vssd1 vccd1 vccd1 _2066_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2753__A _2753_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3849__A _3897_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2175__D _3317_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4390__D _4390_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2968_ _3276_/B _4220_/Q _3150_/S vssd1 vssd1 vccd1 vccd1 _3664_/C sky130_fd_sc_hd__mux2_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2899__S _2941_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1919_ _1941_/A _1918_/Y _4076_/Q vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2899_ _3858_/C _4034_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _3245_/B sky130_fd_sc_hd__mux2_4
XANTENNA__3584__A _3584_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2139__A2 _3879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2928__A _2943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__A _2958_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2075__A1 _4350_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2085__D _2085_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2614__A3 _2421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input88_A gpio_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__C _3925_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2535__C1 _4375_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_5_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output244_A _3160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2550__A2 _2283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2838__A _2898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4120__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2557__B _2557_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4270__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3669__A _3798_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2066__A1 _1952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3940_ _3940_/A _3942_/B _3940_/C vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__and3_1
XANTENNA__2605__A3 _2514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3871_ _3871_/A _3877_/B _3871_/C vssd1 vssd1 vccd1 vccd1 _3872_/A sky130_fd_sc_hd__or3_1
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2822_ _3213_/C _4091_/Q _2858_/S vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__mux2_2
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2753_ _2753_/A vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2369__A2 _2366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1917__A _4356_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2684_ _3283_/B _4118_/Q _3161_/A vssd1 vssd1 vccd1 vccd1 _3457_/C sky130_fd_sc_hd__mux2_1
XFILLER_98_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4354_ _4391_/CLK _4354_/D vssd1 vssd1 vccd1 vccd1 _4354_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2748__A _2748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2541__A2 _3617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3305_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3308_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4285_ _4380_/CLK _4285_/D vssd1 vssd1 vccd1 vccd1 _4285_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4385__D _4385_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3236_ _3250_/A _3236_/B _3250_/C _3245_/D vssd1 vssd1 vccd1 vccd1 _3237_/A sky130_fd_sc_hd__or4_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3167_ _3192_/A _3167_/B _3167_/C _3945_/A vssd1 vssd1 vccd1 vccd1 _3168_/A sky130_fd_sc_hd__and4_1
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2186__C _2186_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _2237_/A _2393_/A _2117_/X vssd1 vssd1 vccd1 vccd1 _2450_/A sky130_fd_sc_hd__a21oi_4
X_3098_ _3227_/C _4201_/Q _3112_/S vssd1 vssd1 vccd1 vccd1 _3620_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3579__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2049_ _2152_/A _3925_/B _3925_/C vssd1 vssd1 vccd1 vccd1 _2050_/D sky130_fd_sc_hd__nand3_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2086__B1_N _4146_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3557__A1 _3557_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3962__D1 _3963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4143__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2532__A2 _4164_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3480__C _4002_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input142_A spi_rty_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4293__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4295__D _4295_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3489__A _3489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2393__A _2393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2599__A2 _2420_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3548__B2 _2530_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3548__A1 _4164_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output194_A _3027_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3655__C _3655_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3952__A _3991_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3671__B _3796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2523__A2 _2362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _4074_/CLK _4070_/D vssd1 vssd1 vccd1 vccd1 _4070_/Q sky130_fd_sc_hd__dfxtp_1
X_3021_ _3021_/A _4242_/Q vssd1 vssd1 vccd1 vccd1 _3022_/A sky130_fd_sc_hd__and2_1
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3484__B1 _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3399__A _3399_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3787__A1 _2117_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3787__B2 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4016__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3923_ _4343_/Q _3908_/A _2024_/Y _3909_/X _3903_/X vssd1 vssd1 vccd1 vccd1 _4343_/D
+ sky130_fd_sc_hd__o2111a_1
X_3854_ _3854_/A vssd1 vssd1 vccd1 vccd1 _4312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2805_ _3204_/B _4088_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _3383_/C sky130_fd_sc_hd__mux2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2750__B _4144_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4166__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3785_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3938_/D sky130_fd_sc_hd__clkbuf_8
X_2736_ _2736_/A vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2667_ _3273_/C _4115_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3451_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3862__A _3862_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2598_ _2319_/X _2248_/X _4172_/Q vssd1 vssd1 vccd1 vccd1 _2598_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3073__S _3073_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4337_ _4356_/CLK _4337_/D vssd1 vssd1 vccd1 vccd1 _4337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4268_ _4282_/CLK _4268_/D vssd1 vssd1 vccd1 vccd1 _4268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2278__A1 _3522_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3219_ _3224_/A _3219_/B _3224_/C _3219_/D vssd1 vssd1 vccd1 vccd1 _3220_/A sky130_fd_sc_hd__or4_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _4199_/CLK _4199_/D vssd1 vssd1 vccd1 vccd1 _4199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__C _2644_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3778__A1 _4276_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3778__B2 input91/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2202__A1 _1930_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3772__A _3772_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2505__A2 _2503_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2593__B1_N _4171_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2483__B_N _2383_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4039__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3012__A _3023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output207_A _2989_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2441__A1 _2439_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3947__A _3976_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4189__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3570_ _3570_/A vssd1 vssd1 vccd1 vccd1 _4181_/D sky130_fd_sc_hd__clkbuf_1
X_2521_ _2519_/Y _2366_/X _2520_/Y vssd1 vssd1 vccd1 vccd1 _2521_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3682__A _3682_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2452_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__buf_4
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2383_ _2383_/A vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2298__A _2298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4172_/CLK _4122_/D vssd1 vssd1 vccd1 vccd1 _4122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4053_ _4074_/CLK _4053_/D vssd1 vssd1 vccd1 vccd1 _4053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3004_ _3010_/A _4234_/Q vssd1 vssd1 vccd1 vccd1 _3005_/A sky130_fd_sc_hd__and2_1
XANTENNA__1930__A _1951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 cpu_adr_i[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2417__D1 _2416_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3279__D _3286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2761__A _2767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3857__A _3881_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3906_ _1987_/Y _3902_/X _1988_/Y _3349_/X _3938_/A vssd1 vssd1 vccd1 vccd1 _4334_/D
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__3576__B _3586_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__A1 _2419_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3837_ _3837_/A _3845_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__and3_1
X_3768_ _4270_/Q _3767_/X _3754_/X input84/X _3755_/X vssd1 vssd1 vccd1 vccd1 _4270_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3295__C _3295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _2719_/A vssd1 vssd1 vccd1 vccd1 _2719_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3932__A1 _2121_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3699_ _3699_/A _4235_/Q _3703_/C _3711_/D vssd1 vssd1 vccd1 vccd1 _3700_/A sky130_fd_sc_hd__and4_1
XANTENNA__3592__A _3804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3160__A2 _2200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2001__A _2001_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2671__A1 _4116_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4331__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A gpio_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3767__A _3767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3486__B _4129_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3923__A1 _4343_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input70_A cpu_sel_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output157_A _2570_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3007__A _3007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2111__B1 _4180_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3677__A _3677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2581__A _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _1952_/A vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3396__B _3405_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3622_ _3635_/A _3635_/B _3622_/C vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__or3_1
XANTENNA__2178__B1 _2177_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3553_ _3553_/A1 _3365_/B _3544_/X _2565_/Y _3547_/X vssd1 vssd1 vccd1 vccd1 _4168_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__1925__A _2022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3484_ _4128_/Q _3350_/X _4395_/A _3469_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _4128_/D
+ sky130_fd_sc_hd__a221o_1
X_2504_ _2287_/X _2424_/X _4162_/Q vssd1 vssd1 vccd1 vccd1 _2504_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__3843__C _3843_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4204__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2435_ _2375_/X _2376_/X _2377_/X _2434_/X _4367_/Q vssd1 vssd1 vccd1 vccd1 _2435_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2350__B1 _2590_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2366_ _2366_/A vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__buf_4
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4105_ _4286_/CLK _4105_/D vssd1 vssd1 vccd1 vccd1 _4105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2297_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2298_/A sky130_fd_sc_hd__buf_4
XANTENNA__4354__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4380_/CLK _4036_/D vssd1 vssd1 vccd1 vccd1 _4036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2503__A_N _2382_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3587__A _3587_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2491__A _4265_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2405__A1 _2379_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2956__A2 _2133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2169__B1 _2013_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput170 _2341_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput192 _3022_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput181 _3000_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2341__B1 _3960_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2666__A _3197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2892__A1 _4033_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3497__A _3497_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4227__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output274_A _2691_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2580__B1 _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4377__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _2517_/A vssd1 vssd1 vccd1 vccd1 _2429_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3960__A _3960_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2332__B1 _2331_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2151_ _2121_/A _3953_/B _4351_/Q vssd1 vssd1 vccd1 vccd1 _2153_/B sky130_fd_sc_hd__o21ai_1
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2082_ _4351_/Q _2182_/B _2081_/Y _1977_/A vssd1 vssd1 vccd1 vccd1 _2083_/D sky130_fd_sc_hd__o211ai_2
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2096__C1 _4250_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2635__A1 _2635_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2984_ _2972_/X _2974_/X _3675_/A vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2399__B1 _2397_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1935_ _2059_/A vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3200__A _3200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3348__C1 _3315_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput50 cpu_dat_i[23] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_2
X_3605_ _3605_/A _3609_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3606_/A sky130_fd_sc_hd__and3_1
Xinput72 cpu_we_i vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_2
Xinput61 cpu_dat_i[4] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 gpio_dat_i[28] vssd1 vssd1 vccd1 vccd1 _2623_/D sky130_fd_sc_hd__clkbuf_2
X_3536_ _3536_/A vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 gpio_dat_i[18] vssd1 vssd1 vccd1 vccd1 _2540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4388__D _4388_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3467_ _3467_/A vssd1 vssd1 vccd1 vccd1 _4121_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3870__A _3870_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2323__B1 _2298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3398_ _3407_/A _3413_/B _3398_/C vssd1 vssd1 vccd1 vccd1 _3399_/A sky130_fd_sc_hd__or3_1
X_2418_ _2418_/A vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2486__A _4264_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2349_ _2349_/A vssd1 vssd1 vccd1 vccd1 _3295_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2917__C _3429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4019_ _4051_/CLK _4019_/D vssd1 vssd1 vccd1 vccd1 _4019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2626__A1 _3560_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2933__B _3447_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3110__A _3117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3051__A1 _4188_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2157__A3 _2153_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2562__B1 _2303_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4298__D _4298_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2396__A _3137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2865__A1 _4098_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input33_A cpu_adr_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3004__B _4234_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2617__B2 _2615_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2617__A1 _2380_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3020__A _3020_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3955__A _3992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4370_ _4380_/CLK _4370_/D vssd1 vssd1 vccd1 vccd1 _4370_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3345__A2 _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2553__B1 _2324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3321_ _3321_/A vssd1 vssd1 vccd1 vccd1 _4062_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3690__A _3690_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3252_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3273_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2305__B1 _2303_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2203_ _2201_/X _1961_/A _1918_/Y _2202_/Y vssd1 vssd1 vccd1 vccd1 _3914_/A sky130_fd_sc_hd__o31ai_4
X_3183_ _3264_/A vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2134_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2662_/A sky130_fd_sc_hd__buf_2
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2456__D _2456_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2065_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2967_ _2197_/X _2200_/X _3661_/A vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3865__A _3865_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2898_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2941_/S sky130_fd_sc_hd__buf_2
X_1918_ _4357_/Q _1923_/A _1924_/A vssd1 vssd1 vccd1 vccd1 _1918_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3584__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3076__S _3076_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3741__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3519_ _3730_/A _2428_/A _3800_/A vssd1 vssd1 vccd1 vccd1 _3547_/A sky130_fd_sc_hd__o21ai_4
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2928__B _2928_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2944__A _2944_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4072__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2075__A2 _2012_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2480__C1 _2469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3925__D _3925_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2535__B1 _2429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2550__A3 _2286_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3015__A _3021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output237_A _3064_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2557__C _2590_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2854__A _2957_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3669__B _3673_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2066__A2 _2160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2605__A4 _2445_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _4319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3685__A _3707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2821_ _3826_/A _4021_/Q _2845_/S vssd1 vssd1 vccd1 vccd1 _3213_/C sky130_fd_sc_hd__mux2_2
X_2752_ _2752_/A _4145_/Q vssd1 vssd1 vccd1 vccd1 _2753_/A sky130_fd_sc_hd__and2_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3971__C1 _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2683_ _2683_/A vssd1 vssd1 vccd1 vccd1 _3161_/A sky130_fd_sc_hd__buf_2
XFILLER_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3723__C1 _3470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4353_ _4391_/CLK _4353_/D vssd1 vssd1 vccd1 vccd1 _4353_/Q sky130_fd_sc_hd__dfxtp_1
X_4284_ _4284_/CLK _4284_/D vssd1 vssd1 vccd1 vccd1 _4284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3304_ _3304_/A vssd1 vssd1 vccd1 vccd1 _4056_/D sky130_fd_sc_hd__clkbuf_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2748__B _4143_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _3235_/A vssd1 vssd1 vccd1 vccd1 _4029_/D sky130_fd_sc_hd__clkbuf_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3707_/A vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__buf_4
XANTENNA__4095__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3097_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _4284_/Q vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__buf_4
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2186__D _2186_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _2182_/A _2081_/B _2053_/A _2081_/D vssd1 vssd1 vccd1 vccd1 _3925_/C sky130_fd_sc_hd__nand4b_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3999_ _3999_/A _3999_/B _4002_/C vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__and3_1
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3557__A2 _3365_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3595__A _3595_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3962__C1 _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2004__A _3294_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2939__A _2939_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input135_A spi_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2599__A3 _2421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3548__A2 _3447_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2756__A0 _4291_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output187_A _2967_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2508__B1 _2507_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3671__C _3675_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3020_ _3020_/A vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3484__A1 _4128_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3484__B2 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3787__A2 _3586_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3922_ _2167_/Y _3902_/X _2013_/Y _3566_/A _3331_/X vssd1 vssd1 vccd1 vccd1 _4342_/D
+ sky130_fd_sc_hd__o2111ai_1
X_3853_ _3871_/A _3853_/B _3853_/C vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__or3_1
XFILLER_60_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2804_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2851_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__1928__A input7/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3784_ _4282_/Q _3657_/A _3771_/A input98/X _3772_/A vssd1 vssd1 vccd1 vccd1 _4282_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2735_ _2737_/A _4137_/Q vssd1 vssd1 vccd1 vccd1 _2736_/A sky130_fd_sc_hd__and2_1
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2666_ _3197_/A vssd1 vssd1 vccd1 vccd1 _2947_/S sky130_fd_sc_hd__buf_2
XANTENNA__2759__A _3197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2597_ _2592_/X _2596_/Y _2499_/X _2579_/X vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__o211a_1
X_4336_ _4356_/CLK _4336_/D vssd1 vssd1 vccd1 vccd1 _4336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _4286_/CLK _4267_/D vssd1 vssd1 vccd1 vccd1 _4267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2278__A2 _2255_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4198_ _4275_/CLK _4198_/D vssd1 vssd1 vccd1 vccd1 _4198_/Q sky130_fd_sc_hd__dfxtp_1
X_3218_ _3218_/A vssd1 vssd1 vccd1 vccd1 _4023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3149_ _3149_/A vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3778__A2 _3767_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_4_CLK_A clkbuf_2_1_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2435__C1 _4367_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4110__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2202__A2 _2201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4260__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2910__A0 _3863_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2441__A2 _3673_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2520_ _2575_/A _2520_/B _2520_/C _2520_/D vssd1 vssd1 vccd1 vccd1 _2520_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__3963__A _3963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2451_ _2363_/X _2449_/X _2311_/X _2450_/X _4368_/Q vssd1 vssd1 vccd1 vccd1 _2451_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2579__A _2579_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3154__B1 _3569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2382_ _2382_/A vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _4251_/CLK _4121_/D vssd1 vssd1 vccd1 vccd1 _4121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4052_ _4085_/CLK _4052_/D vssd1 vssd1 vccd1 vccd1 _4052_/Q sky130_fd_sc_hd__dfxtp_1
X_3003_ _3003_/A vssd1 vssd1 vccd1 vccd1 _3003_/X sky130_fd_sc_hd__clkbuf_1
Xinput4 cpu_adr_i[11] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3203__A _3343_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4133__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2417__C1 _2409_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2968__A0 _3276_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3905_ _3940_/C vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2761__B _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__A2 _3535_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3576__C _3576_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3836_ _3884_/A vssd1 vssd1 vccd1 vccd1 _3855_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3767_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3767_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4283__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2718_ _2726_/A _4129_/Q vssd1 vssd1 vccd1 vccd1 _2719_/A sky130_fd_sc_hd__and2_1
XANTENNA__3873__A _3897_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3932__A2 _2201_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3698_ _4234_/Q _3695_/X _3696_/X _3697_/X _3683_/X vssd1 vssd1 vccd1 vccd1 _4234_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2649_ _2328_/A _2329_/A _2469_/A _2648_/Y vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4371_/CLK _4319_/D vssd1 vssd1 vccd1 vccd1 _4319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3113__A _3117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2959__A0 _3180_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3486__C _3502_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3923__A2 _3908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2592__D1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input63_A cpu_dat_i[6] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3023__A _3023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4156__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output317_A _2194_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2111__A1 _2087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__C1 _4389_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3958__A _3958_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1952_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3396__C _3400_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3621_ _3621_/A vssd1 vssd1 vccd1 vccd1 _4201_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3693__A _3699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3552_ _3558_/A _3552_/B vssd1 vssd1 vccd1 vccd1 _4167_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2178__A1 _4067_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2503_ _2382_/X _2383_/X _2503_/C _2503_/D vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__1925__B _2023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3483_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2102__A _2638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2434_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__buf_2
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2365_ _4257_/Q vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _4180_/CLK _4104_/D vssd1 vssd1 vccd1 vccd1 _4104_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2350__A1 _4250_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1941__A _1941_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2296_ _2367_/A _2393_/A _2336_/A vssd1 vssd1 vccd1 vccd1 _2533_/A sky130_fd_sc_hd__and3_1
XFILLER_57_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4035_ _4199_/CLK _4035_/D vssd1 vssd1 vccd1 vccd1 _4035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3868__A _3868_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2405__A2 _2399_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3819_ _3823_/A _3829_/B _3819_/C vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__or3_1
XANTENNA__2169__A1 _2167_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4029__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3108__A _3127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput160 _2597_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2012__A _2167_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput182 _3003_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[15] sky130_fd_sc_hd__buf_2
Xoutput193 _3025_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[25] sky130_fd_sc_hd__buf_2
XFILLER_88_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput171 _2359_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__4179__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2341__A1 _2328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2385__C _2385_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output267_A _2747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3109__A0 _3236_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3018__A _3018_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2580__A1 _2512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__B _3973_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2332__A1 _2332_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2150_ _2150_/A _2182_/B vssd1 vssd1 vccd1 vccd1 _2153_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2081_ _2150_/A _2081_/B _2081_/C _2081_/D vssd1 vssd1 vccd1 vccd1 _2081_/Y sky130_fd_sc_hd__nand4b_2
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2096__B1 _4286_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2635__A2 _2628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2983_ _3291_/C _4225_/Q _3157_/S vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2399__B2 _2398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2399__A1 _2380_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1934_ _1934_/A vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3348__B1 _2063_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput40 cpu_dat_i[14] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1936__A _3916_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput73 gpio_ack_i vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
Xinput51 cpu_dat_i[24] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3604_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3624_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput62 cpu_dat_i[5] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
Xinput95 gpio_dat_i[29] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_2
Xinput84 gpio_dat_i[19] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_2
X_3535_ _3546_/A _3535_/B vssd1 vssd1 vccd1 vccd1 _4155_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4004__B1_N _2648_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2571__A1 _2423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3466_ _3466_/A _3584_/B _3466_/C vssd1 vssd1 vccd1 vccd1 _3467_/A sky130_fd_sc_hd__and3_1
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4321__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2417_ _2406_/X _2407_/X _2408_/X _2409_/X _2416_/Y vssd1 vssd1 vccd1 vccd1 _2417_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2767__A _2767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2323__A1 _4254_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3397_ _3397_/A vssd1 vssd1 vccd1 vccd1 _4093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2323__B2 input99/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2348_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2406_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2279_ _2224_/X _2245_/X _2246_/X _3949_/A vssd1 vssd1 vccd1 vccd1 _2279_/X sky130_fd_sc_hd__o211a_2
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4085_/CLK _4018_/D vssd1 vssd1 vccd1 vccd1 _4018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2626__A2 _2526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3598__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2933__C _3437_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3110__B _3125_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2007__A _2007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2562__A1 _2427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2562__B2 _2304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2677__A _2752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2484__B1_N _4160_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2396__B _3677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A cpu_adr_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2617__A2 _2614_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3301__A _3301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4344__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2437__B1_N _4156_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2553__B2 _2552_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2553__A1 _2301_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3320_ _3320_/A _3320_/B _3326_/C _3326_/D vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__or4_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2305__A1 _2301_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3251_ _3251_/A vssd1 vssd1 vccd1 vccd1 _4036_/D sky130_fd_sc_hd__clkbuf_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2305__B2 _2304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3182_ _3953_/C vssd1 vssd1 vccd1 vccd1 _3264_/A sky130_fd_sc_hd__buf_2
X_2202_ _1930_/X _2201_/A _1994_/X _4337_/Q vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__o31ai_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _2133_/A vssd1 vssd1 vccd1 vccd1 _2133_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2064_ _4075_/Q _2152_/A _2063_/Y vssd1 vssd1 vccd1 vccd1 _2064_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2069__B1 _2068_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3211__A _3211_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2966_ _3273_/C _4219_/Q _3335_/A vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3865__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2241__B1 _2113_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2897_ _4314_/Q input50/X _2940_/S vssd1 vssd1 vccd1 vccd1 _3858_/C sky130_fd_sc_hd__mux2_1
X_1917_ _4356_/Q vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__inv_2
XANTENNA__3584__C _3600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2544__A1 _2386_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3741__B1 _2315_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3881__A _3881_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3518_ _2225_/Y _3308_/A _3469_/X _3470_/A vssd1 vssd1 vccd1 vccd1 _4146_/D sky130_fd_sc_hd__a211oi_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3449_ _3457_/A _3462_/B _3449_/C vssd1 vssd1 vccd1 vccd1 _3450_/A sky130_fd_sc_hd__or3_1
XANTENNA__3092__S _3112_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2928__C _3434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4217__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2480__B1 _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4367__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3980__B1 _2494_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1991__C1 _1990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4102__D _4102_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2535__B2 _2434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2535__A1 _2481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3791__A _3884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2200__A _2200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2299__B1 _2298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3015__B _4239_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2557__D _2557_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3669__C _3669_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3031__A _3031_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2870__A _3197_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2820_ _4301_/Q input36/X _2844_/S vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__mux2_8
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _2751_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3971__B1 _2442_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2682_ _3891_/C _4048_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _3283_/B sky130_fd_sc_hd__mux2_4
XFILLER_99_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4012__D _4012_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__B1 _3044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4352_ _4391_/CLK _4352_/D vssd1 vssd1 vccd1 vccd1 _4352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4283_ _4284_/CLK _4283_/D vssd1 vssd1 vccd1 vccd1 _4283_/Q sky130_fd_sc_hd__dfxtp_1
X_3303_ _3320_/A _3303_/B _3317_/C _3326_/D vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__or4_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3206__A _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3234_ _3247_/A _3253_/B _3234_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _3235_/A sky130_fd_sc_hd__and4_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ _3953_/C vssd1 vssd1 vccd1 vccd1 _3707_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2116_ input73/X _2272_/A _2272_/B _2115_/Y vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__o31a_4
X_3096_ _3099_/A _3106_/B _3618_/C vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__and3_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2047_ _2120_/A _2141_/A _4345_/Q vssd1 vssd1 vccd1 vccd1 _3925_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__2483__C _2483_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3876__A _3876_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2780__A _2799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3998_ _3991_/X _3992_/X _2617_/Y vssd1 vssd1 vccd1 vccd1 _4385_/D sky130_fd_sc_hd__o21bai_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3557__A3 _3544_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2214__B1 _2213_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2949_ _4288_/Q input68/X _2949_/S vssd1 vssd1 vccd1 vccd1 _3794_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3962__B1 _2357_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2004__B _3294_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2020__A _2020_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input128_A spi_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input93_A gpio_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2205__B1 _1949_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2756__A1 input35/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2508__A1 _2506_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3026__A _3032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3484__A2 _3350_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2692__A0 _4330_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3696__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3921_ _4341_/Q _3908_/X _2028_/Y _3909_/X _3903_/X vssd1 vssd1 vccd1 vccd1 _4341_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3852_ _3876_/A vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4007__D _4007_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2803_ _3819_/C _4018_/Q _2826_/S vssd1 vssd1 vccd1 vccd1 _3204_/B sky130_fd_sc_hd__mux2_4
XANTENNA__1928__B _1970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3783_ _3769_/A _3764_/A _3748_/A _2639_/Y _3774_/X vssd1 vssd1 vccd1 vccd1 _4281_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3944__B1 _3728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2105__A _4391_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2734_ _2734_/A vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__clkbuf_1
X_2665_ _2683_/A vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1944__A _1951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2596_ _2526_/X _3556_/B _2595_/Y vssd1 vssd1 vccd1 vccd1 _2596_/Y sky130_fd_sc_hd__o21ai_2
X_4335_ _4356_/CLK _4335_/D vssd1 vssd1 vccd1 vccd1 _4335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4062__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2253__B1_N _4147_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4266_ _4280_/CLK _4266_/D vssd1 vssd1 vccd1 vccd1 _4266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4197_ _4275_/CLK _4197_/D vssd1 vssd1 vccd1 vccd1 _4197_/Q sky130_fd_sc_hd__dfxtp_1
X_3217_ _3221_/A _3227_/B _3217_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__and4_1
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2775__A _2896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _3151_/A _3657_/B _3653_/A vssd1 vssd1 vccd1 vccd1 _3149_/A sky130_fd_sc_hd__and3_1
XFILLER_83_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3079_ _3115_/A vssd1 vssd1 vccd1 vccd1 _3109_/S sky130_fd_sc_hd__buf_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2435__B1 _2377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2015__A _2055_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2202__A3 _1994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4392__318 vssd1 vssd1 vccd1 vccd1 _4392__318/HI cpu_err_o sky130_fd_sc_hd__conb_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2371__C1 _2370_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2910__A1 _4036_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2674__A0 _3889_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2426__B1 _2425_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output297_A _2913_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4085__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3963__B _3973_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2450_ _2450_/A vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__buf_4
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3154__A1 _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2381_ _2543_/A vssd1 vssd1 vccd1 vccd1 _3536_/A sky130_fd_sc_hd__clkbuf_2
X_4120_ _4250_/CLK _4120_/D vssd1 vssd1 vccd1 vccd1 _4120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4051_/CLK _4051_/D vssd1 vssd1 vccd1 vccd1 _4051_/Q sky130_fd_sc_hd__dfxtp_1
X_3002_ _3010_/A _4233_/Q vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__and2_1
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 cpu_adr_i[12] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2417__B1 _2408_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2968__A1 _4220_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3904_ input33/X _3902_/X _2002_/Y _3938_/D _3903_/X vssd1 vssd1 vccd1 vccd1 _4333_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__1939__A input8/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2761__C _3367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3835_ _3835_/A vssd1 vssd1 vccd1 vccd1 _4304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3766_ _3752_/X _3764_/X _3765_/X _2541_/Y _3757_/X vssd1 vssd1 vccd1 vccd1 _4269_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3917__B1 _1946_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2717_ _2739_/A vssd1 vssd1 vccd1 vccd1 _2726_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3932__A3 _1994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3697_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2648_ _2526_/X _2645_/Y _2509_/X _2646_/Y _2647_/Y vssd1 vssd1 vccd1 vccd1 _2648_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4200__D _4200_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2579_ _2579_/A vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4391_/CLK _4318_/D vssd1 vssd1 vccd1 vccd1 _4318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4249_ _4282_/CLK _4249_/D vssd1 vssd1 vccd1 vccd1 _4249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3113__B _3125_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2959__A1 _4080_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2592__C1 _2409_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input56_A cpu_dat_i[29] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4110__D _4110_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3304__A _3304_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2111__A2 _2226_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__B1 _2429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output212_A _3087_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _2059_/A vssd1 vssd1 vccd1 vccd1 _1962_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3974__A _3974_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3620_ _3620_/A _3633_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__and3_1
XANTENNA__3693__B _4233_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3551_ _3551_/A1 _3536_/X _3544_/X _2549_/Y _3537_/X vssd1 vssd1 vccd1 vccd1 _4166_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__2178__A2 _2093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2502_ _2481_/X _2501_/X _2377_/X _2434_/X _4373_/Q vssd1 vssd1 vccd1 vccd1 _2502_/X
+ sky130_fd_sc_hd__o221a_1
X_3482_ _3876_/A vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__buf_6
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2433_ _2417_/X _2432_/Y _2404_/X _2373_/X vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__o211a_2
XANTENNA_clkbuf_leaf_3_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2364_ _2363_/X _2258_/X _2311_/X _2260_/X _4364_/Q vssd1 vssd1 vccd1 vccd1 _2364_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2886__A0 _3853_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__D _4020_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2350__A2 _3295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4103_ _4275_/CLK _4103_/D vssd1 vssd1 vccd1 vccd1 _4103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2295_ _3720_/A vssd1 vssd1 vccd1 vccd1 _2295_/X sky130_fd_sc_hd__buf_4
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4100__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3214__A _3214_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4034_ _4380_/CLK _4034_/D vssd1 vssd1 vccd1 vccd1 _4034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4250__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3884__A _3884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3818_ _3818_/A vssd1 vssd1 vccd1 vccd1 _4297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2169__A2 _3902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3095__S _3109_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3749_ _3727_/X _3747_/X _3748_/X _2416_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _4259_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput161 _2603_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput150 _2511_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__2012__B _2012_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput194 _3027_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput183 _3005_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2877__A0 _3236_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2326__C1 _2325_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput172 _2374_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__2341__A2 _2329_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2629__B1 _2628_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2385__D _2503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input110_A spi_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4105__D _4105_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3794__A _3798_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3109__A1 _4204_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output162_A _2612_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2580__A2 _2513_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4123__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2317__C1 _2316_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__C _3963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2868__A0 _4309_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2332__A2 _2090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3034__A _3036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4273__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2080_ _2204_/A _2018_/X _4071_/Q vssd1 vssd1 vccd1 vccd1 _2083_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__2873__A _2873_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3969__A _3992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2096__A1 _1965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2635__A3 _2514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2982_ _2972_/X _2974_/X _3673_/C vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2399__A2 _2389_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ _1930_/X _1932_/X _4338_/Q vssd1 vssd1 vccd1 vccd1 _3916_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__4015__D _4015_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3603_ _3603_/A vssd1 vssd1 vccd1 vccd1 _4194_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3348__A1 _4075_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput30 cpu_adr_i[6] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_2
XANTENNA__1936__B _3916_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput52 cpu_dat_i[25] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_2
Xinput41 cpu_dat_i[15] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3209__A _3209_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput63 cpu_dat_i[6] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
Xinput96 gpio_dat_i[2] vssd1 vssd1 vccd1 vccd1 _2314_/D sky130_fd_sc_hd__clkbuf_1
Xinput85 gpio_dat_i[1] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_2
Xinput74 gpio_dat_i[0] vssd1 vssd1 vccd1 vccd1 _2275_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3534_ _3549_/A vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2113__A _2113_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2571__A2 _2446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3465_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3584_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2416_ _2410_/Y _2411_/X _2415_/Y vssd1 vssd1 vccd1 vccd1 _2416_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__1952__A _1952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2767__B _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2323__A2 _2322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3396_ _3396_/A _3405_/B _3400_/C vssd1 vssd1 vccd1 vccd1 _3397_/A sky130_fd_sc_hd__and3_1
XFILLER_97_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2347_ _3730_/A vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__buf_6
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2278_ _3522_/B _2255_/X _2261_/Y _2277_/Y vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__o211ai_4
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2783__A _3447_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3879__A _3879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4017_ _4051_/CLK _4017_/D vssd1 vssd1 vccd1 vccd1 _4017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3598__B _3611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3110__C _3626_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3119__A _3137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4146__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2023__A _2023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2562__A2 _2428_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4296__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2396__C _2507_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A cpu_adr_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3301__B _3328_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3029__A _3029_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2002__A1 _1930_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2553__A2 _2302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3250_/A _3250_/B _3250_/C _3271_/D vssd1 vssd1 vccd1 vccd1 _3251_/A sky130_fd_sc_hd__or4_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2305__A2 _2302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3181_ _3181_/A vssd1 vssd1 vccd1 vccd1 _4010_/D sky130_fd_sc_hd__clkbuf_1
X_2201_ _2201_/A vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__clkbuf_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _3343_/B vssd1 vssd1 vccd1 vccd1 _2133_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__A _3699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2069__A1 _2134_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2063_ _2061_/Y _2001_/A _2062_/Y _2059_/A vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4019__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2108__A _2113_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4169__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2965_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3335_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2241__A1 _4286_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2896_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2940_/S sky130_fd_sc_hd__buf_2
XANTENNA__3865__C _3879_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2544__B1_N _4165_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3517_ _3517_/A vssd1 vssd1 vccd1 vccd1 _4145_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2544__A2 _2424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3741__A1 _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3448_ _3448_/A vssd1 vssd1 vccd1 vccd1 _4113_/D sky130_fd_sc_hd__clkbuf_1
X_3379_ _3379_/A vssd1 vssd1 vccd1 vccd1 _4086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3402__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2480__A1 _2328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2018__A _2018_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2232__A1 _2422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3980__A1 _3968_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__B2 _2498_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1991__B1 _1986_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2535__A2 _2501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2688__A _2898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2299__A1 _4252_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2299__B2 input85/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__A _3332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2471__A1 _2330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4311__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2750_ _2752_/A _4144_/Q vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__and2_1
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3971__A1 _4367_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2681_ _4328_/Q input28/X _2949_/S vssd1 vssd1 vccd1 vccd1 _3891_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3982__A _3982_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__A1 _4248_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__B2 _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4351_ _4356_/CLK _4351_/D vssd1 vssd1 vccd1 vccd1 _4351_/Q sky130_fd_sc_hd__dfxtp_1
X_4282_ _4282_/CLK _4282_/D vssd1 vssd1 vccd1 vccd1 _4282_/Q sky130_fd_sc_hd__dfxtp_1
X_3302_ _3302_/A vssd1 vssd1 vccd1 vccd1 _4055_/D sky130_fd_sc_hd__clkbuf_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3233_ _3692_/A vssd1 vssd1 vccd1 vccd1 _3253_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ input1/X vssd1 vssd1 vccd1 vccd1 _3953_/C sky130_fd_sc_hd__buf_2
X_3095_ _3224_/B _4200_/Q _3109_/S vssd1 vssd1 vccd1 vccd1 _3618_/C sky130_fd_sc_hd__mux2_1
X_2115_ _4284_/Q vssd1 vssd1 vccd1 vccd1 _2115_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3222__A _3222_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2046_ _2204_/A _2018_/A _4065_/Q vssd1 vssd1 vccd1 vccd1 _2050_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__2483__D _2503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2780__B _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3997_ _3997_/A vssd1 vssd1 vccd1 vccd1 _4384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2948_ _2677_/X _2680_/X _3354_/A vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2214__A1 _2139_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3962__A1 _2342_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2879_ _2879_/A vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4203__D _4203_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3892__A _3892_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2004__C _2145_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2301__A _2427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3132__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4334__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2205__A1 _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input86_A gpio_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4113__D _4113_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2610__D1 _2609_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2910__S _2941_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2508__A2 _2411_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3307__A _3433_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2211__A _2211_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3026__B _4244_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output242_A _3156_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2692__A1 input30/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3042__A _3120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3977__A _3977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3920_ _2006_/Y _3902_/X _2008_/Y _3349_/X _3331_/X vssd1 vssd1 vccd1 vccd1 _4340_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3851_ _3851_/A vssd1 vssd1 vccd1 vccd1 _4311_/D sky130_fd_sc_hd__clkbuf_1
X_3782_ _4280_/Q _3657_/A _3771_/X input95/X _3772_/X vssd1 vssd1 vccd1 vccd1 _4280_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3929__D1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2802_ _4298_/Q input64/X _2825_/S vssd1 vssd1 vccd1 vccd1 _3819_/C sky130_fd_sc_hd__mux2_2
X_2733_ _2737_/A _4136_/Q vssd1 vssd1 vccd1 vccd1 _2734_/A sky130_fd_sc_hd__and2_1
XANTENNA__3944__A1 _2407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3944__B2 _2552_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4023__D _4023_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2820__S _2844_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4207__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2664_ _3885_/A _4045_/Q _2936_/S vssd1 vssd1 vccd1 vccd1 _3273_/C sky130_fd_sc_hd__mux2_2
X_2595_ _2301_/X _2428_/X _2303_/X _2304_/X _4382_/Q vssd1 vssd1 vccd1 vccd1 _2595_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3217__A _3221_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2121__A _2121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4334_ _4347_/CLK _4334_/D vssd1 vssd1 vccd1 vccd1 _4334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4286_/CLK _4265_/D vssd1 vssd1 vccd1 vccd1 _4265_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4357__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1960__A _2078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4196_ _4275_/CLK _4196_/D vssd1 vssd1 vccd1 vccd1 _4196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3216_ _3216_/A vssd1 vssd1 vccd1 vccd1 _4022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147_ _3265_/C _4215_/Q _3147_/S vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3078_ _3078_/A vssd1 vssd1 vccd1 vccd1 _3078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3887__A _3895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2435__B2 _2434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2435__A1 _2375_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2029_ _4341_/Q _1970_/A _2028_/Y _2015_/X _2136_/A vssd1 vssd1 vccd1 vccd1 _2030_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3098__S _3112_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1946__B1 _4339_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3127__A _3127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2031__A _2031_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2360__B1_N _4153_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2371__B1 _2364_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input140_A spi_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2123__B1 _3945_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2674__A1 _4047_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2186__A_N _3326_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4108__D _4108_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3797__A _3797_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2426__A1 _2426_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2905__S _2905_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output192_A _3022_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1937__B1 _1936_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__C _3963_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3154__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3037__A _3037_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2380_ _2380_/A vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__buf_4
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4050_ _4326_/CLK _4050_/D vssd1 vssd1 vccd1 vccd1 _4050_/Q sky130_fd_sc_hd__dfxtp_1
X_3001_ _3023_/A vssd1 vssd1 vccd1 vccd1 _3010_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2114__B1 _3945_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 cpu_adr_i[13] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4018__D _4018_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3500__A _3500_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2417__A1 _2406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2815__S _2825_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__clkbuf_2
X_3834_ _3847_/A _3853_/B _3834_/C vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__or3_1
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3917__A1 _1939_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3765_ _3765_/A vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1955__A _4357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__clkbuf_2
X_2716_ _2716_/A vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__clkbuf_1
Xoutput310 _2813_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[8] sky130_fd_sc_hd__buf_2
X_2647_ _2427_/X _2501_/X _2429_/X _2430_/X _4389_/Q vssd1 vssd1 vccd1 vccd1 _2647_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2578_ _3554_/B _2362_/X _2573_/Y _2577_/Y vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__o211ai_4
X_4317_ _4371_/CLK _4317_/D vssd1 vssd1 vccd1 vccd1 _4317_/Q sky130_fd_sc_hd__dfxtp_1
X_4248_ _4264_/CLK _4248_/D vssd1 vssd1 vccd1 vccd1 _4248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4179_ _4180_/CLK _4179_/D vssd1 vssd1 vccd1 vccd1 _4179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3113__C _3629_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__A _3410_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1919__B1 _4076_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2592__B1 _2408_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input49_A cpu_dat_i[22] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2647__A1 _2427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__B2 _2430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output205_A _2984_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3320__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3693__C _3703_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3550_ _3558_/A _3550_/B vssd1 vssd1 vccd1 vccd1 _4165_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3780__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2501_ _3730_/B vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__clkbuf_4
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _4127_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3990__A _3990_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4301__D _4301_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2432_ _2419_/X _3535_/B _2431_/Y vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2363_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__buf_4
XANTENNA__2886__A1 _4032_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _4180_/CLK _4102_/D vssd1 vssd1 vccd1 vccd1 _4102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2294_ _3578_/A vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4033_ _4199_/CLK _4033_/D vssd1 vssd1 vccd1 vccd1 _4033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3230__A _3295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3817_ _3817_/A _3821_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__and3_1
X_3748_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3748_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3679_ _4226_/Q _3351_/X _4394_/A _3678_/X _3504_/X vssd1 vssd1 vccd1 vccd1 _4226_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4211__D _4211_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2326__B1 _2293_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput151 _2525_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput195 _3029_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput184 _3007_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[17] sky130_fd_sc_hd__buf_2
Xoutput162 _2612_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_82_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2877__A1 _4100_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput173 _2405_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_88_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3405__A _3405_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2629__B2 _2286_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2629__A1 _3466_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4075__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3140__A _3140_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input103_A gpio_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3794__B _3805_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3762__C1 _3757_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__D _4121_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2317__B1 _2312_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2868__A1 input44/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2332__A3 _2308_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3315__A _3315_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output155_A _2307_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3034__B _4248_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2096__A2 _1942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2635__A4 _2531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3050__A _3050_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _3288_/B _4224_/Q _3150_/S vssd1 vssd1 vccd1 vccd1 _3673_/C sky130_fd_sc_hd__mux2_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ _2007_/A vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__buf_2
Xinput20 cpu_adr_i[26] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
X_3602_ _3611_/A _3611_/B _3602_/C vssd1 vssd1 vccd1 vccd1 _3603_/A sky130_fd_sc_hd__or3_1
XANTENNA__3348__A2 _3314_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput31 cpu_adr_i[7] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1936__C _1977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput53 cpu_dat_i[26] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_0_CLK_A CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput42 cpu_dat_i[16] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput64 cpu_dat_i[7] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_4
Xinput97 gpio_dat_i[30] vssd1 vssd1 vccd1 vccd1 _2638_/D sky130_fd_sc_hd__buf_2
Xinput86 gpio_dat_i[20] vssd1 vssd1 vccd1 vccd1 _2557_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 gpio_dat_i[10] vssd1 vssd1 vccd1 vccd1 _2456_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3533_ _2385_/C _3523_/X _3528_/X _2388_/Y _3562_/A vssd1 vssd1 vccd1 vccd1 _4154_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3753__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__D _4031_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3464_ _3800_/A vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__buf_2
XFILLER_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3505__C1 _3504_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2415_ _2507_/A _2557_/B _2590_/C _2415_/D vssd1 vssd1 vccd1 vccd1 _2415_/Y sky130_fd_sc_hd__nand4_1
XFILLER_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2767__C _3370_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3395_ _3395_/A vssd1 vssd1 vccd1 vccd1 _4092_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3225__A _3225_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4098__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2346_ _2346_/A vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__buf_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2277_ _2262_/X _2375_/A _2408_/A _2409_/A _2276_/Y vssd1 vssd1 vccd1 vccd1 _2277_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_4016_ _4085_/CLK _4016_/D vssd1 vssd1 vccd1 vccd1 _4016_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3879__B _3893_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3598__C _3598_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3895__A _3895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__D _4206_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2795__A0 _4297_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2304__A _2552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2547__B1 _2546_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3744__C1 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3135__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2396__D _2396_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2180__D1 _2136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2974__A _3326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3301__C _3695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4116__D _4116_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_2_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2786__A0 _3192_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output272_A _2676_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2002__A2 _1932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4240__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2200_ _2200_/A vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3045__A _3045_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3180_ _3195_/A _3180_/B _3195_/C _3190_/D vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__or4_1
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2884__A _2884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2131_ _2678_/A vssd1 vssd1 vccd1 vccd1 _3343_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3699__B _4235_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4390__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2062_ _1952_/A _2007_/A _4355_/Q vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2069__A2 _3935_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2108__B _2108_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2964_ _2964_/A vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__buf_2
XANTENNA__4026__D _4026_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2895_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2241__A2 _2349_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2124__A _4002_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3726__C1 _3470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3516_ _3516_/A _4145_/Q _3657_/C vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__and3_1
XANTENNA__3741__A2 _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3447_ _3447_/A _3447_/B _4002_/B vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__and3_1
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3378_ _3383_/A _3389_/B _3378_/C vssd1 vssd1 vccd1 vccd1 _3379_/A sky130_fd_sc_hd__or3_1
XFILLER_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2329_ _2329_/A vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2794__A _2957_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2162__D1 _1965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3402__B _3413_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2480__A2 _2329_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4113__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2232__A2 _2446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__A2 _3969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4263__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1991__A1 _1976_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2940__A0 _4322_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2299__A2 _2295_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A cpu_adr_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2604__B1_N _4173_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2471__A2 _2446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2619__B1_N _4175_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3971__A2 _3965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2680_ _3190_/D vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__buf_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2879__A _2879_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3982__B _3999_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4356_/CLK _4350_/D vssd1 vssd1 vccd1 vccd1 _4350_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3723__A2 _3167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2931__A0 _3871_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3301_ _3301_/A _3328_/B _3695_/A _3925_/D vssd1 vssd1 vccd1 vccd1 _3302_/A sky130_fd_sc_hd__and4_1
XFILLER_99_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4281_ _4286_/CLK _4281_/D vssd1 vssd1 vccd1 vccd1 _4281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3232_ _3232_/A vssd1 vssd1 vccd1 vccd1 _4028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3163_ _3335_/A vssd1 vssd1 vccd1 vccd1 _3167_/B sky130_fd_sc_hd__buf_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3503__A _3503_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2114_ _4286_/Q _2349_/A _3945_/D vssd1 vssd1 vccd1 vccd1 _2517_/A sky130_fd_sc_hd__o21ai_4
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3094_ _3094_/A vssd1 vssd1 vccd1 vccd1 _3094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4136__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2045_ _4344_/Q _1970_/A _2044_/Y _1938_/A vssd1 vssd1 vccd1 vccd1 _2050_/B sky130_fd_sc_hd__o211ai_1
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1958__A _2078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2780__C _3374_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3996_ _3996_/A _3999_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__and3_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2214__A2 _3115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4286__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2947_ _3167_/C _4077_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3354_/A sky130_fd_sc_hd__mux2_2
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3962__A2 _2357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2878_ _2888_/A _2901_/B _3413_/C vssd1 vssd1 vccd1 vccd1 _2879_/A sky130_fd_sc_hd__and3_1
XANTENNA__2004__D _2145_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2922__A0 _3257_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3413__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3132__B _3142_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2205__A2 _1996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2610__C1 _2454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input79_A gpio_dat_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4009__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2211__B _2211_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output235_A _3058_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4159__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3323__A _3343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3977__B _3999_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3850_ _3850_/A _3869_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__and3_1
X_2801_ _3489_/A vssd1 vssd1 vccd1 vccd1 _2828_/A sky130_fd_sc_hd__clkbuf_1
X_3781_ _3769_/X _3764_/A _3748_/A _2624_/Y _3774_/X vssd1 vssd1 vccd1 vccd1 _4279_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3929__C1 _3909_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2732_ _2732_/A vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2601__C1 _4383_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3944__A2 _2406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4304__D _4304_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3157__A0 _3178_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2663_ _2958_/S vssd1 vssd1 vccd1 vccd1 _2936_/S sky130_fd_sc_hd__buf_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2594_ _2594_/A1 _3369_/A _2286_/A _2593_/Y vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__a31oi_4
XANTENNA__2904__A0 _4315_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3217__B _3227_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4333_ _4347_/CLK _4333_/D vssd1 vssd1 vccd1 vccd1 _4333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4264_ _4264_/CLK _4264_/D vssd1 vssd1 vccd1 vccd1 _4264_/Q sky130_fd_sc_hd__dfxtp_1
X_3215_ _3224_/A _3215_/B _3224_/C _3219_/D vssd1 vssd1 vccd1 vccd1 _3216_/A sky130_fd_sc_hd__or4_1
XFILLER_68_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4195_ _4199_/CLK _4195_/D vssd1 vssd1 vccd1 vccd1 _4195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3233__A _3692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3146_ _3146_/A vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3077_ _3081_/A _3089_/B _3605_/A vssd1 vssd1 vccd1 vccd1 _3078_/A sky130_fd_sc_hd__and3_1
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2071__A2_N _4070_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ _2028_/A _2072_/B _2081_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2028_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3887__B _3935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2435__A2 _2376_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4214__D _4214_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3979_ _4371_/Q _3965_/X _2489_/Y _3966_/Y vssd1 vssd1 vccd1 vccd1 _4371_/D sky130_fd_sc_hd__a211o_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1946__A1 _2120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3408__A _3408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2031__B _3320_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2371__A1 _3532_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4301__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3143__A _3143_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2123__A1 _4391_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input133_A spi_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2426__A2 _2420_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4124__D _4124_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2921__S _2941_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1937__A1 _4058_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output185_A _3009_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3318__A _3318_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3053__A _3053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2114__A1 _4286_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3000_ _3000_/A vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__clkbuf_1
Xinput7 cpu_adr_i[14] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2417__A2 _2407_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3902_ _3902_/A vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__clkbuf_2
X_3833_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3853_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4034__D _4034_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2831__S _2844_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3917__A2 _3902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2715_ _2715_/A _4128_/Q vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__and2_1
X_3695_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1955__B _2201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput300 _2929_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[28] sky130_fd_sc_hd__buf_2
X_2646_ _4282_/Q _2295_/X _2298_/X input98/X vssd1 vssd1 vccd1 vccd1 _2646_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__2132__A _3343_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3228__A _3228_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1998__A_N input32/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4324__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput311 _2819_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2577_ _2474_/X _2452_/X _2453_/X _2454_/X _2576_/Y vssd1 vssd1 vccd1 vccd1 _2577_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _4391_/CLK _4316_/D vssd1 vssd1 vccd1 vccd1 _4316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _4282_/CLK _4247_/D vssd1 vssd1 vccd1 vccd1 _4247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4178_ _4388_/CLK _4178_/D vssd1 vssd1 vccd1 vccd1 _4178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4209__D _4209_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3898__A _3898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3129_ _3135_/A _3142_/B _3638_/A vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__and3_1
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__B _3429_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1919__A1 _1941_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2577__D1 _2576_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2041__B1 _2040_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2592__A1 _2376_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2977__A _3115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2647__A2 _2501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4119__D _4119_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3_0_CLK_A clkbuf_2_3_0_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2916__S _2916_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3601__A _3601_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__B _3320_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__D1 _3938_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4347__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3693__D _3711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3480_ _3492_/A _4127_/Q _4002_/B vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__and3_1
XANTENNA__3780__B1 _3771_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2500_ _2494_/X _2498_/Y _2499_/X _2469_/X vssd1 vssd1 vccd1 vccd1 _2500_/X sky130_fd_sc_hd__o211a_1
X_2431_ _2427_/X _2428_/X _2429_/X _2430_/X _4366_/Q vssd1 vssd1 vccd1 vccd1 _2431_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2362_ _2380_/A vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__buf_4
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2293_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2293_/X sky130_fd_sc_hd__buf_4
X_4101_ _4275_/CLK _4101_/D vssd1 vssd1 vccd1 vccd1 _4101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4032_ _4380_/CLK _4032_/D vssd1 vssd1 vccd1 vccd1 _4032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4029__D _4029_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3511__A _3511_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2826__S _2826_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2127__A _2700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3816_ _3816_/A vssd1 vssd1 vccd1 vccd1 _4296_/D sky130_fd_sc_hd__clkbuf_1
X_3747_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2559__D1 _2558_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__clkbuf_2
X_2629_ _3466_/C _4176_/Q _2628_/X _2286_/X vssd1 vssd1 vccd1 vccd1 _2629_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_82_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2326__A1 _2281_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput152 _2537_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput185 _3009_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput163 _2618_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[27] sky130_fd_sc_hd__buf_2
XANTENNA__2326__B2 _2323_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput174 _2433_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[8] sky130_fd_sc_hd__buf_2
Xoutput196 _3031_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[28] sky130_fd_sc_hd__buf_2
XANTENNA__3405__B _3405_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2629__A2 _4176_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3421__A _3421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2037__A _2037_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3794__C _3794_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2565__A1 _2319_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3762__B1 _2521_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input61_A cpu_dat_i[4] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2317__A1 _3527_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2332__A4 _2421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output148_A _2490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output315_A _2960_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2096__A3 _1918_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3331__A _3940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _2972_/X _2974_/X _3671_/A vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1931_ _4356_/Q _2023_/A _2022_/A vssd1 vssd1 vccd1 vccd1 _2007_/A sky130_fd_sc_hd__nand3b_2
Xinput21 cpu_adr_i[27] vssd1 vssd1 vccd1 vccd1 _2150_/A sky130_fd_sc_hd__buf_2
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _4193_/D sky130_fd_sc_hd__clkbuf_1
Xinput10 cpu_adr_i[17] vssd1 vssd1 vccd1 vccd1 _2027_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 cpu_dat_i[27] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_2
XANTENNA__3753__B1 _2457_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4312__D _4312_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput43 cpu_dat_i[17] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 cpu_adr_i[8] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 gpio_dat_i[21] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
Xinput98 gpio_dat_i[31] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_2
Xinput76 gpio_dat_i[11] vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__clkbuf_1
X_3532_ _3564_/B _3532_/B vssd1 vssd1 vccd1 vccd1 _4153_/D sky130_fd_sc_hd__nor2_1
Xinput65 cpu_dat_i[8] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
X_3463_ _3463_/A vssd1 vssd1 vccd1 vccd1 _4120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3505__B1 _3489_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3506__A _3976_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2414_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2590_/C sky130_fd_sc_hd__buf_2
XANTENNA__2410__A _4259_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3394_ _3407_/A _3413_/B _3394_/C vssd1 vssd1 vccd1 vccd1 _3395_/A sky130_fd_sc_hd__or3_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2345_ _2366_/A vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__buf_2
X_2276_ _2268_/Y _2539_/A _2275_/Y vssd1 vssd1 vccd1 vccd1 _2276_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3879__C _3879_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4015_ _4051_/CLK _4015_/D vssd1 vssd1 vccd1 vccd1 _4015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3241__A _3250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3895__B _3935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2795__A1 input63/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4222__D _4222_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3744__B1 _3735_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2547__A1 _2419_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3416__A _3416_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_21_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4199_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3135__B _3142_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4042__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2180__C1 _1973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4192__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3151__A _3151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2990__A _3036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3301__D _3925_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2786__A1 _4085_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4132__D _4132_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output265_A _2743_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3326__A _3343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4284_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2130_ _2130_/A vssd1 vssd1 vccd1 vccd1 _2678_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3699__C _3703_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2061_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3061__A _3061_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3996__A _3996_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4307__D _4307_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ _2197_/X _2200_/X _3659_/C vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2894_ _2917_/A _2901_/B _3420_/A vssd1 vssd1 vccd1 vccd1 _2895_/A sky130_fd_sc_hd__and3_1
XANTENNA__4042__D _4042_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3726__B1 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3515_ _4144_/Q _3308_/A _2767_/A _3490_/A _3504_/X vssd1 vssd1 vccd1 vccd1 _4144_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4065__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__A3 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3236__A _3250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3446_ _3976_/A vssd1 vssd1 vccd1 vccd1 _4002_/B sky130_fd_sc_hd__buf_2
XFILLER_100_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3377_ _3377_/A vssd1 vssd1 vccd1 vccd1 _4085_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2162__C1 _1973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2328_ _2328_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2259_ _2517_/A vssd1 vssd1 vccd1 vccd1 _3728_/A sky130_fd_sc_hd__buf_4
XFILLER_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3402__C _3402_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4217__D _4217_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2217__B1 _3052_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1991__A2 _1977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3146__A _3146_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A1 input59/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2050__A _2050_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2985__A _3023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input24_A cpu_adr_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4127__D _4127_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4371_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2225__A _2700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4088__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3982__C _3996_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2931__A1 _4040_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3300_ _3300_/A vssd1 vssd1 vccd1 vccd1 _4054_/D sky130_fd_sc_hd__clkbuf_1
X_4280_ _4280_/CLK _4280_/D vssd1 vssd1 vccd1 vccd1 _4280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2895__A _2895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3231_ _3250_/A _3231_/B _3250_/C _3245_/D vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__or4_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3192_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2144__C1 _3303_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2695__B1 _3462_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2113_ _2113_/A vssd1 vssd1 vccd1 vccd1 _3945_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3099_/A _3106_/B _3614_/A vssd1 vssd1 vccd1 vccd1 _3094_/A sky130_fd_sc_hd__and3_1
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2044_ _2044_/A _2081_/B _2053_/A _2081_/D vssd1 vssd1 vccd1 vccd1 _2044_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__4037__D _4037_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3995_ _3991_/X _3992_/X _2602_/Y vssd1 vssd1 vccd1 vccd1 _4383_/D sky130_fd_sc_hd__o21bai_1
X_2946_ _3792_/A _4007_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _3167_/C sky130_fd_sc_hd__mux2_1
X_2877_ _3236_/B _4100_/Q _2911_/S vssd1 vssd1 vccd1 vccd1 _3413_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2922__A1 _4108_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3429_ _3429_/A _3429_/B _3455_/C vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_1_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__B _3413_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2438__B1 _2437_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3132__C _3642_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4230__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2610__B1 _2453_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4380__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2374__C1 _2373_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2211__C _2211_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3604__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3323__B _3326_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output228_A _3140_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3977__C _3996_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2800_ _2800_/A vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__clkbuf_1
X_3780_ _4278_/Q _3767_/X _3771_/X input93/X _3772_/X vssd1 vssd1 vccd1 vccd1 _4278_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3929__B1 _2038_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2731_ _2737_/A _4135_/Q vssd1 vssd1 vccd1 vccd1 _2732_/A sky130_fd_sc_hd__and2_1
XANTENNA__2601__B1 _2324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3157__A1 _4183_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2662_ _2662_/A vssd1 vssd1 vccd1 vccd1 _2958_/S sky130_fd_sc_hd__buf_2
X_2593_ _2386_/X _2289_/X _4171_/Q vssd1 vssd1 vccd1 vccd1 _2593_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__4320__D _4320_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2904__A1 input51/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3217__C _3217_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4332_ _4356_/CLK _4332_/D vssd1 vssd1 vccd1 vccd1 _4332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4263_ _4286_/CLK _4263_/D vssd1 vssd1 vccd1 vccd1 _4263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3514__A _3514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4103__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3214_ _3214_/A vssd1 vssd1 vccd1 vccd1 _4021_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2668__B1 _3451_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4194_ _4286_/CLK _4194_/D vssd1 vssd1 vccd1 vccd1 _4194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _3151_/A _3657_/B _3650_/C vssd1 vssd1 vccd1 vccd1 _3146_/A sky130_fd_sc_hd__and3_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4253__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3076_ _3213_/C _4195_/Q _3076_/S vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__mux2_2
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2027_ _2027_/A vssd1 vssd1 vccd1 vccd1 _2028_/A sky130_fd_sc_hd__inv_2
XANTENNA__1969__A _2093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3887__C _3887_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2840__A0 _3219_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A vssd1 vssd1 vccd1 vccd1 _4370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2929_ _2929_/A vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1946__A2 _2141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4230__D _4230_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2031__C _2031_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2371__A2 _2362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3424__A _3424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2123__A2 _2357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input126_A spi_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2426__A3 _2421_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2831__A0 _4303_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input91_A gpio_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2595__C1 _4382_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1937__A2 _2184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output178_A _2994_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__D _4140_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4276__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2114__A2 _2349_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput8 cpu_adr_i[15] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2822__A0 _3213_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3901_ _3900_/X _1998_/Y _3470_/X _3314_/X vssd1 vssd1 vccd1 vccd1 _4332_/D sky130_fd_sc_hd__a211o_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4315__D _4315_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3832_ _3832_/A vssd1 vssd1 vccd1 vccd1 _4303_/D sky130_fd_sc_hd__clkbuf_1
X_3763_ _4268_/Q _3750_/X _3754_/X input82/X _3755_/X vssd1 vssd1 vccd1 vccd1 _4268_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2586__C1 _4381_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2714_ _2714_/A vssd1 vssd1 vccd1 vccd1 _2714_/X sky130_fd_sc_hd__clkbuf_1
X_3694_ _3694_/A vssd1 vssd1 vccd1 vccd1 _4233_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2413__A _2590_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput301 _2934_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[29] sky130_fd_sc_hd__buf_2
X_2645_ _3444_/A _4178_/Q _2644_/X _2286_/X vssd1 vssd1 vccd1 vccd1 _2645_/Y sky130_fd_sc_hd__a22oi_2
Xoutput312 _2948_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__4050__D _4050_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2576_ _2574_/Y _2366_/X _2575_/Y vssd1 vssd1 vccd1 vccd1 _2576_/Y sky130_fd_sc_hd__o21ai_4
X_4315_ _4371_/CLK _4315_/D vssd1 vssd1 vccd1 vccd1 _4315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1971__B _1998_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3244__A _3244_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4246_ _4264_/CLK _4246_/D vssd1 vssd1 vccd1 vccd1 _4246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4177_/CLK _4177_/D vssd1 vssd1 vccd1 vccd1 _4177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3128_ _3247_/C _4209_/Q _3147_/S vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3898__B _3942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3195_/B _4190_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3594_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3066__A0 _3204_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3410__C _3424_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4225__D _4225_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4149__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3419__A _3419_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2577__C1 _2454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1919__A2 _1918_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2041__A1 _2036_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2592__A2 _2375_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4299__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2993__A _2999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__C _3326_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4135__D _4135_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2932__S _2942_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4006__C1 _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output295_A _2902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2568__C1 _4379_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3329__A _3329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3780__A1 _4278_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3780__B2 input93/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2430_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3064__A _3064_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2361_ _2361_/A1 _2090_/A _2308_/X _2421_/A _2360_/Y vssd1 vssd1 vccd1 vccd1 _3532_/B
+ sky130_fd_sc_hd__a41oi_4
X_4100_ _4180_/CLK _4100_/D vssd1 vssd1 vccd1 vccd1 _4100_/Q sky130_fd_sc_hd__dfxtp_1
X_2292_ _2292_/A vssd1 vssd1 vccd1 vccd1 _2509_/A sky130_fd_sc_hd__buf_2
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3999__A _3999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4031_ _4199_/CLK _4031_/D vssd1 vssd1 vccd1 vccd1 _4031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3296__B1 _3346_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2408__A _2408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3048__A0 _3188_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4001__B1_N _2632_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4045__D _4045_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3815_ _3823_/A _3829_/B _3815_/C vssd1 vssd1 vccd1 vccd1 _3816_/A sky130_fd_sc_hd__or3_1
X_3746_ _4258_/Q _3734_/X _3735_/X _2396_/D _3738_/X vssd1 vssd1 vccd1 vccd1 _4258_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2559__C1 _2409_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3239__A _3247_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3677_ _3677_/A vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__buf_2
XANTENNA__1982__A _2078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2628_ _2628_/A _2644_/B _2628_/C vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__and3_1
XANTENNA__2326__A2 _2321_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput186 _3011_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput164 _2627_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2559_ _2406_/X _2375_/X _2408_/X _2409_/X _2558_/Y vssd1 vssd1 vccd1 vccd1 _2559_/X
+ sky130_fd_sc_hd__o2111a_2
Xoutput153 _2548_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput175 _2443_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput197 _3033_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[29] sky130_fd_sc_hd__buf_2
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3405__C _3424_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _4262_/CLK _4229_/D vssd1 vssd1 vccd1 vccd1 _4229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3702__A _3720_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3039__A0 _3184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3149__A _3149_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2053__A _2053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2565__A2 _2289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3762__A1 _3752_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2988__A _2988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input54_A cpu_dat_i[27] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2317__A2 _2255_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2927__S _2937_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3612__A _3612_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output210_A _3078_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output308_A _2800_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4314__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2253__A1 _2644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 cpu_adr_i[28] vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__clkbuf_2
X_3600_ _3600_/A _3609_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__and3_1
Xinput11 cpu_adr_i[18] vssd1 vssd1 vccd1 vccd1 _2167_/A sky130_fd_sc_hd__buf_2
Xinput55 cpu_dat_i[28] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3753__A1 _3752_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3531_ _2353_/Y _3523_/X _2356_/A _3349_/X _2419_/X vssd1 vssd1 vccd1 vccd1 _4152_/D
+ sky130_fd_sc_hd__o2111ai_1
Xinput44 cpu_dat_i[18] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput33 cpu_adr_i[9] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_2
Xinput88 gpio_dat_i[22] vssd1 vssd1 vccd1 vccd1 _2575_/D sky130_fd_sc_hd__clkbuf_2
Xinput77 gpio_dat_i[12] vssd1 vssd1 vccd1 vccd1 _2476_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2898__A _2898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput66 cpu_dat_i[9] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_2
Xinput99 gpio_dat_i[3] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_2
X_3462_ _3586_/A _3462_/B _3462_/C vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__or3_1
XANTENNA__3505__A1 _4138_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3505__B2 _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3393_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3413_/B sky130_fd_sc_hd__clkbuf_2
X_2413_ _2590_/B vssd1 vssd1 vccd1 vccd1 _2557_/B sky130_fd_sc_hd__buf_2
X_2344_ _2344_/A vssd1 vssd1 vccd1 vccd1 _2366_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3910__D1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3522__A _3564_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2275_ _2412_/A _2590_/B _2414_/A _2275_/D vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__2837__S _2885_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4014_ _4085_/CLK _4014_/D vssd1 vssd1 vccd1 vccd1 _4014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3241__B _3241_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1977__A _1977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3895__C _3895_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3744__A1 _4256_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2547__A2 _3550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3744__B2 _3744_/B2 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3729_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3135__C _3644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2180__B1 _2179_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3432__A _3432_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4337__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3151__B _3657_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2640__D1 _2639_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3607__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output160_A _2597_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3326__B _3326_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output258_A _2668_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2657__S _2942_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__D _3711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2060_ _4073_/Q _2152_/A _2059_/Y vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3996__B _3999_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2962_ _3271_/B _4218_/Q _3150_/S vssd1 vssd1 vccd1 vccd1 _3659_/C sky130_fd_sc_hd__mux2_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2388__B1_N _4154_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2893_ _3243_/C _4103_/Q _2916_/S vssd1 vssd1 vccd1 vccd1 _3420_/A sky130_fd_sc_hd__mux2_4
XANTENNA__4323__D _4323_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3726__A1 _2099_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3514_ _3514_/A vssd1 vssd1 vccd1 vccd1 _4143_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3517__A _3517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2421__A _2421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3445_ _3953_/C vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3236__B _3236_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3376_ _3376_/A _3381_/B _3376_/C vssd1 vssd1 vccd1 vccd1 _3377_/A sky130_fd_sc_hd__and3_1
XANTENNA__2162__B1 _2161_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2224_/X _2245_/X _2326_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__o211a_2
XANTENNA__3252__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2258_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__buf_4
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2189_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2864_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2217__A1 _2197_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4233__D _4233_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3427__A _3427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2050__B _2050_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3162__A _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A cpu_adr_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2506__A _4266_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3956__A1 _3952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4143__D _4143_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2940__S _2940_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3337__A _3800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _3295_/C vssd1 vssd1 vccd1 vccd1 _3250_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__2144__B1 _1990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2695__A1 _2677_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _3161_/A vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__buf_4
XANTENNA__3341__C1 _3346_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A _3127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2112_ _2129_/B _2112_/B vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _3221_/C _4199_/Q _3112_/S vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4318__D _4318_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2447__A1 _2330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3800__A _3800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2043_ _2043_/A vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__inv_2
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _3968_/X _3969_/X _2592_/X _2596_/Y vssd1 vssd1 vccd1 vccd1 _4382_/D sky130_fd_sc_hd__o22a_1
XANTENNA__4032__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4053__D _4053_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2945_ _4287_/Q input67/X _2953_/S vssd1 vssd1 vccd1 vccd1 _3792_/A sky130_fd_sc_hd__mux2_1
X_2876_ _3847_/C _4030_/Q _2886_/S vssd1 vssd1 vccd1 vccd1 _3236_/B sky130_fd_sc_hd__mux2_4
XANTENNA__2850__S _2886_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4182__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3247__A _3247_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3428_ _3428_/A vssd1 vssd1 vccd1 vccd1 _3455_/C sky130_fd_sc_hd__buf_2
XANTENNA__2135__A0 _4323_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3359_ _3359_/A vssd1 vssd1 vccd1 vccd1 _4078_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input9_A cpu_adr_i[16] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3413__C _3413_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4228__D _4228_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2438__A1 _3536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2610__A1 _2474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2760__S _2955_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2061__A _2061_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2374__B1 _3963_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2996__A _2996_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2211__D _2211_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3323__C _3323_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4138__D _4138_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3620__A _3620_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2935__S _2935_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4055__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3929__A1 _4347_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2730_ _2730_/A vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2601__B2 _2552_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2601__A1 _2407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2670__S _2950_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2661_ _4325_/Q input13/X _2935_/S vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__mux2_8
XANTENNA__3067__A _3081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2592_ _2376_/X _2375_/X _2408_/X _2409_/X _2591_/Y vssd1 vssd1 vccd1 vccd1 _2592_/X
+ sky130_fd_sc_hd__o2111a_2
XANTENNA__3217__D _3234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4331_ _4346_/CLK _4331_/D vssd1 vssd1 vccd1 vccd1 _4331_/Q sky130_fd_sc_hd__dfxtp_1
X_4262_ _4262_/CLK _4262_/D vssd1 vssd1 vccd1 vccd1 _4262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3213_ _3221_/A _3227_/B _3213_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _3214_/A sky130_fd_sc_hd__and4_1
XANTENNA__2668__A1 _2128_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4199_/CLK _4193_/D vssd1 vssd1 vccd1 vccd1 _4193_/Q sky130_fd_sc_hd__dfxtp_1
X_3144_ _3262_/B _4214_/Q _3144_/S vssd1 vssd1 vccd1 vccd1 _3650_/C sky130_fd_sc_hd__mux2_1
X_3075_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2845__S _2845_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4048__D _4048_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3530__A _3564_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2026_ _2204_/A _2018_/X _4061_/Q vssd1 vssd1 vccd1 vccd1 _2030_/C sky130_fd_sc_hd__o21ai_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2840__A1 _4094_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2146__A _2146_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3977_ _3977_/A _3999_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__and3_1
XANTENNA__1985__A _2055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _2943_/A _2928_/B _3434_/A vssd1 vssd1 vccd1 vccd1 _2929_/A sky130_fd_sc_hd__and3_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2859_/A _2872_/B _3405_/A vssd1 vssd1 vccd1 vccd1 _2860_/A sky130_fd_sc_hd__and3_1
XANTENNA__3553__C1 _3547_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3705__A _3935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3424__B _3429_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4078__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3440__A _3440_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input119_A spi_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2831__A1 input38/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input84_A gpio_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2595__B1 _2303_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3615__A _3615_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output240_A _3075_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 cpu_adr_i[16] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3350__A _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2822__A1 _4091_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _1971_/C _1971_/D _1998_/B _4332_/Q vssd1 vssd1 vccd1 vccd1 _3900_/X sky130_fd_sc_hd__a31o_1
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3831_ _3831_/A _3845_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__and3_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3762_ _3752_/X _3747_/X _3748_/X _2521_/Y _3757_/X vssd1 vssd1 vccd1 vccd1 _4267_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_0_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__C1 _3774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2586__B1 _2429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2713_ _2715_/A _4127_/Q vssd1 vssd1 vccd1 vccd1 _2714_/A sky130_fd_sc_hd__and2_1
X_3693_ _3699_/A _4233_/Q _3703_/C _3711_/D vssd1 vssd1 vccd1 vccd1 _3694_/A sky130_fd_sc_hd__and4_1
XANTENNA__4331__D _4331_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2644_ _2644_/A _2644_/B _2644_/C vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__and3_1
Xoutput302 _2774_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput313 _2952_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[1] sky130_fd_sc_hd__buf_2
X_2575_ _2575_/A _2638_/B _2638_/C _2575_/D vssd1 vssd1 vccd1 vccd1 _2575_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__2338__B1 _2337_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3525__A _3547_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4314_ _4380_/CLK _4314_/D vssd1 vssd1 vccd1 vccd1 _4314_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1971__C _1971_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4220__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4245_ _4282_/CLK _4245_/D vssd1 vssd1 vccd1 vccd1 _4245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _4389_/CLK _4176_/D vssd1 vssd1 vccd1 vccd1 _4176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3127_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3142_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2510__B1 _2508_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3898__C _3914_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4370__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3260__A _3273_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3058_ _3058_/A vssd1 vssd1 vccd1 vccd1 _3058_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3066__A1 _4192_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ _2006_/Y _2168_/A _2008_/Y _2137_/A _1985_/X vssd1 vssd1 vccd1 vccd1 _2009_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2577__B1 _2453_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4241__D _4241_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2041__A2 _1962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3526__C1 _3562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3435__A _3435_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2993__B _4229_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3170__A _3201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__D _3326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4006__B1 _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2514__A _2514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2568__B1 _2324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output190_A _3018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output288_A _2867_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4151__D _4151_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3780__A2 _3767_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4243__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2360_ _2330_/X _2424_/A _4153_/Q vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2291_ _3526_/A1 _2283_/X _2286_/X _2290_/Y vssd1 vssd1 vccd1 vccd1 _2291_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3999__B _3999_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4030_ _4380_/CLK _4030_/D vssd1 vssd1 vccd1 vccd1 _4030_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3296__A1 _2145_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3048__A1 _4187_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4326__D _4326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2424__A _2424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2559__B1 _2408_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _4295_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3756__C1 _3755_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3745_ _3727_/X _3729_/X _3732_/X _2369_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _4257_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3239__B _3253_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4061__D _4061_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3676_ _3676_/A vssd1 vssd1 vccd1 vccd1 _4225_/D sky130_fd_sc_hd__clkbuf_1
X_2627_ _2581_/X _2582_/X _3999_/A _2246_/X vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3255__A _3297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput143 _2125_/X vssd1 vssd1 vccd1 vccd1 cpu_ack_o sky130_fd_sc_hd__buf_2
Xoutput176 _2963_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput165 _2633_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_88_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2558_ _2556_/Y _3617_/A _2557_/Y vssd1 vssd1 vccd1 vccd1 _2558_/Y sky130_fd_sc_hd__o21ai_4
Xoutput154 _2555_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput198 _2969_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[2] sky130_fd_sc_hd__buf_2
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput187 _2967_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[1] sky130_fd_sc_hd__buf_2
X_2489_ _2380_/X _2485_/Y _2488_/X _2398_/X vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2072__A_N input18/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4228_ _4262_/CLK _4228_/D vssd1 vssd1 vccd1 vccd1 _4228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4159_ _4180_/CLK _4159_/D vssd1 vssd1 vccd1 vccd1 _4159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3039__A1 _4185_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4116__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4236__D _4236_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2798__A0 _3199_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2334__A _4255_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4266__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2053__B _2074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3762__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2988__B _4227_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2970__A0 _3279_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3165__A _3953_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input47_A cpu_dat_i[20] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2509__A _2509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4146__D _4146_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output203_A _2980_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2789__A0 _4296_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2253__A2 _2424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2244__A _2582_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 cpu_adr_i[19] vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 cpu_adr_i[29] vssd1 vssd1 vccd1 vccd1 _2057_/C sky130_fd_sc_hd__buf_2
X_3530_ _3564_/B _3530_/B vssd1 vssd1 vccd1 vccd1 _4151_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3753__A2 _3747_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput45 cpu_dat_i[19] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 cpu_cyc_i vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__clkbuf_4
Xinput89 gpio_dat_i[23] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_2
Xinput78 gpio_dat_i[13] vssd1 vssd1 vccd1 vccd1 _2487_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 cpu_dat_i[29] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_2
Xinput67 cpu_sel_i[0] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_4
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3075__A _3075_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3505__A2 _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2412_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2507_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3392_ _3392_/A vssd1 vssd1 vccd1 vccd1 _4091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2343_ _4256_/Q vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3910__C1 _3909_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3803__A _3803_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3522__B _3522_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2274_ _2638_/C vssd1 vssd1 vccd1 vccd1 _2414_/A sky130_fd_sc_hd__clkbuf_2
X_4013_ _4051_/CLK _4013_/D vssd1 vssd1 vccd1 vccd1 _4013_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4139__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2419__A _2526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3241__C _3250_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4056__D _4056_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4289__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3744__A2 _3734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1993__A _2204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1989_ _1987_/Y _2168_/A _1988_/Y _1977_/A vssd1 vssd1 vccd1 vccd1 _1989_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__2952__B1 _3358_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3728_ _3728_/A vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__buf_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3659_ _3659_/A _3659_/B _3659_/C vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__or3_1
XANTENNA__3901__C1 _3314_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2180__A1 _2044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2329__A _2329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3151__C _3655_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2048__B _2081_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2763__S _2953_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input101_A gpio_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2640__C1 _2454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2999__A _2999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3607__B _3611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3326__C _3326_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A _3623_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output153_A _2548_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2459__C1 _2458_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__S _2935_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3996__C _3996_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2961_ _3115_/A vssd1 vssd1 vccd1 vccd1 _3150_/S sky130_fd_sc_hd__buf_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2631__C1 _4387_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2892_ _3855_/A _4033_/Q _2905_/S vssd1 vssd1 vccd1 vccd1 _3243_/C sky130_fd_sc_hd__mux2_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2702__A _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3726__A2 _3167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3513_ _3516_/A _4143_/Q _3657_/C vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__and3_1
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3444_ _3444_/A vssd1 vssd1 vccd1 vccd1 _3447_/A sky130_fd_sc_hd__buf_2
XANTENNA__3236__C _3250_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2147__D1 _2069_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3375_ _3375_/A vssd1 vssd1 vccd1 vccd1 _4084_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2162__A1 _2024_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2281_/X _2321_/Y _2293_/X _2323_/Y _2325_/Y vssd1 vssd1 vccd1 vccd1 _2326_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2257_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2474_/A sky130_fd_sc_hd__clkbuf_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2188_ _2188_/A _2211_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__nand3_4
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2217__A2 _2200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2495__B1_N _4161_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3708__A _3717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2925__A0 _4319_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4304__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2050__C _2050_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3443__A _3443_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2758__S _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2059__A _2059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3102__A0 _3231_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3956__A2 _3955_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3618__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2916__A0 _3253_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output270_A _2751_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3353__A _3444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2144__A1 _2140_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _2988_/A _2200_/A _3576_/C vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3341__B1 _3340_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2695__A2 _2680_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3091_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3106_/B sky130_fd_sc_hd__clkbuf_1
X_2111_ _2087_/A _2226_/A _4180_/Q vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__a21oi_4
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2042_ _1993_/X _2018_/X _4064_/Q vssd1 vssd1 vccd1 vccd1 _2050_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2447__A2 _2446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _3991_/X _3992_/X _2587_/Y vssd1 vssd1 vccd1 vccd1 _4381_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__4334__D _4334_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2944_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3528__A _3544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2875_ _4310_/Q input45/X _2885_/S vssd1 vssd1 vccd1 vccd1 _3847_/C sky130_fd_sc_hd__mux2_2
XANTENNA__2080__B1 _4071_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4327__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3247__B _3253_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3427_ _3427_/A vssd1 vssd1 vccd1 vccd1 _4106_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3263__A _3263_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2135__A1 input72/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3358_ _3470_/A _3365_/B _3358_/C vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__or3_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2644_/A _2424_/A _4149_/Q vssd1 vssd1 vccd1 vccd1 _2309_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3289_ _3289_/A vssd1 vssd1 vccd1 vccd1 _4050_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2438__A2 _2436_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2607__A _4277_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4244__D _4244_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2610__A2 _2452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2071__B1 _2015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3438__A _3438_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2342__A _4363_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2374__A1 _2328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3173__A _3343_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2517__A _2517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3112__S _3112_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3620__B _3633_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4154__D _4154_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2951__S _3161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3929__A2 _3908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2601__A2 _2302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2062__B1 _4355_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2252__A _2514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2660_ _2957_/S vssd1 vssd1 vccd1 vccd1 _2935_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3067__B _3070_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2591_ _2589_/Y _3617_/A _2590_/Y vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_5_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4347_/CLK _4330_/D vssd1 vssd1 vccd1 vccd1 _4330_/Q sky130_fd_sc_hd__dfxtp_1
X_4261_ _4286_/CLK _4261_/D vssd1 vssd1 vccd1 vccd1 _4261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3083__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3212_ _3264_/A vssd1 vssd1 vccd1 vccd1 _3234_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2668__A2 _2133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2522__D1 _2521_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4192_ _4286_/CLK _4192_/D vssd1 vssd1 vccd1 vccd1 _4192_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4329__D _4329_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3143_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3811__A _3811_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3074_ _3081_/A _3089_/B _3602_/C vssd1 vssd1 vccd1 vccd1 _3075_/A sky130_fd_sc_hd__and3_1
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3530__B _3530_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2427__A _2427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2025_ _4343_/Q _1970_/A _2024_/Y _2015_/X _1985_/X vssd1 vssd1 vccd1 vccd1 _2030_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_91_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2146__B _2146_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4064__D _4064_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _3999_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2927_ _3260_/C _4109_/Q _2937_/S vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3258__A _3258_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2858_ _3227_/C _4097_/Q _2858_/S vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__mux2_4
X_2789_ _4296_/Q input62/X _2825_/S vssd1 vssd1 vccd1 vccd1 _3815_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3553__B1 _2565_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3424__C _3424_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4239__D _4239_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3721__A _3767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2337__A _2412_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2771__S _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2595__B2 _2304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2595__A1 _2301_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3168__A _3168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2503__C _2503_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input77_A gpio_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2800__A _2800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4149__D _4149_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4022__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output233_A _3152_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3631__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2946__S _2954_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2247__A _2446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4172__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2681__S _2949_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3830_ _3830_/A vssd1 vssd1 vccd1 vccd1 _4302_/D sky130_fd_sc_hd__clkbuf_1
X_3761_ _4266_/Q _3750_/X _3754_/X _2507_/D _3755_/X vssd1 vssd1 vccd1 vccd1 _4266_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2035__B1 _2034_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2712_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3078__A _3078_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2586__A1 _2481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2586__B2 _2430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__B1 _2639_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3692_ _3692_/A vssd1 vssd1 vccd1 vccd1 _3711_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2643_ _3428_/A vssd1 vssd1 vccd1 vccd1 _3444_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2338__A1 _2334_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput303 _2939_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2710__A _2710_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput314 _2956_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[2] sky130_fd_sc_hd__buf_2
X_2574_ _4273_/Q vssd1 vssd1 vccd1 vccd1 _2574_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3806__A _3806_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4313_ _4371_/CLK _4313_/D vssd1 vssd1 vccd1 vccd1 _4313_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1971__D _1971_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _4264_/CLK _4244_/D vssd1 vssd1 vccd1 vccd1 _4244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4175_ _4177_/CLK _4175_/D vssd1 vssd1 vccd1 vccd1 _4175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3541__A _3546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4059__D _4059_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3126_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2510__B2 _2509_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2510__A1 _2255_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3260__B _3279_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3057_ _3063_/A _3070_/B _3589_/A vssd1 vssd1 vccd1 vccd1 _3058_/A sky130_fd_sc_hd__and3_1
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3471__C1 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1996__A _2018_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2008_ _2120_/A _2160_/A _4340_/Q vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2026__B1 _4061_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2577__A1 _2474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3959_ _3952_/X _3955_/X _2326_/Y vssd1 vssd1 vccd1 vccd1 _4361_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__3526__B1 _2290_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4045__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2766__S _2937_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4195__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input131_A spi_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3451__A _3451_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A1 _4391_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2017__B1 _2016_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2568__A1 _2301_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2568__B2 _2552_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output183_A _3005_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2530__A _2628_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3626__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ _2287_/X _2289_/X _4148_/Q vssd1 vssd1 vccd1 vccd1 _2290_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3999__C _4002_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3361__A _3361_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3296__A2 _2145_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2705__A _2705_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2008__B1 _4340_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3813_ _3813_/A _3821_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__and3_1
XANTENNA__2559__A1 _2406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4342__D _4342_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3756__B1 _3754_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3744_ _4256_/Q _3734_/X _3735_/X _3744_/B2 _3738_/X vssd1 vssd1 vccd1 vccd1 _4256_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3239__C _3239_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3675_ _3675_/A _3796_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__and3_1
XANTENNA__3536__A _3536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2440__A _2507_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2626_ _3560_/B _2526_/A _2621_/Y _2625_/Y vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__o211ai_4
Xoutput177 _2992_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2557_ _2590_/A _2557_/B _2590_/C _2557_/D vssd1 vssd1 vccd1 vccd1 _2557_/Y sky130_fd_sc_hd__nand4_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput155 _2307_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput144 _2279_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput166 _2318_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput199 _3035_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[30] sky130_fd_sc_hd__buf_2
Xoutput188 _3014_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[20] sky130_fd_sc_hd__buf_2
X_2488_ _2486_/Y _2411_/X _2487_/Y vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__o21a_4
X_4227_ _4262_/CLK _4227_/D vssd1 vssd1 vccd1 vccd1 _4227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3271__A _3276_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4158_ _4172_/CLK _4158_/D vssd1 vssd1 vccd1 vccd1 _4158_/Q sky130_fd_sc_hd__dfxtp_1
X_3109_ _3236_/B _4204_/Q _3109_/S vssd1 vssd1 vccd1 vccd1 _3626_/C sky130_fd_sc_hd__mux2_1
X_4089_ _4225_/CLK _4089_/D vssd1 vssd1 vccd1 vccd1 _4089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2798__A1 _4087_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4252__D _4252_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2053__C _2053_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3762__A3 _3748_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3446__A _3976_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_2_3_0_CLK clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2970__A1 _4221_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_24_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3181__A _3181_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2385__B_N _2383_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2238__B1 _4283_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2789__A1 input62/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4162__D _4162_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4210__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 cpu_adr_i[1] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
Xinput46 cpu_dat_i[1] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 cpu_dat_i[0] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
Xinput24 cpu_adr_i[2] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_4
Xinput79 gpio_dat_i[14] vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3356__A _3591_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3753__A3 _3748_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2260__A _2552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4360__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput68 cpu_sel_i[1] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_4
Xinput57 cpu_dat_i[2] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_15_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4264_/CLK sky130_fd_sc_hd__clkbuf_16
X_3460_ _3460_/A vssd1 vssd1 vccd1 vccd1 _4119_/D sky130_fd_sc_hd__clkbuf_1
X_2411_ _3641_/A vssd1 vssd1 vccd1 vccd1 _2411_/X sky130_fd_sc_hd__clkbuf_4
X_3391_ _3391_/A _3405_/B _3400_/C vssd1 vssd1 vccd1 vccd1 _3392_/A sky130_fd_sc_hd__and3_1
X_2342_ _4363_/Q vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3910__B1 _1983_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3091__A _3127_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2273_ _2336_/A vssd1 vssd1 vccd1 vccd1 _2638_/C sky130_fd_sc_hd__clkbuf_2
X_4012_ _4051_/CLK _4012_/D vssd1 vssd1 vccd1 vccd1 _4012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2477__B1 _2476_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3241__D _3245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4337__D _4337_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2229__B1 _2356_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4072__D _4072_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3727_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1988_ _1930_/X _2141_/A _4334_/Q vssd1 vssd1 vccd1 vccd1 _1988_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2952__A1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__A _3266_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3658_ _3658_/A vssd1 vssd1 vccd1 vccd1 _4217_/D sky130_fd_sc_hd__clkbuf_1
X_2609_ _2607_/Y _2366_/A _2608_/Y vssd1 vssd1 vccd1 vccd1 _2609_/Y sky130_fd_sc_hd__o21ai_4
X_3589_ _3589_/A _3609_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__and3_1
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3901__B1 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2165__C1 _2184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2180__A2 _2001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__B1 _2467_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4247__D _4247_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2048__C _2053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4233__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2345__A _2366_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2033__B1_N _4346_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2640__B1 _2453_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4383__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2999__B _4232_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3176__A _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3607__C _3607_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3326__D _3326_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output146_A _2470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2459__B1 _2451_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4157__D _4157_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output313_A _2952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2954__S _2954_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4388_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _2704_/A _2133_/A _3365_/C vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2255__A _2418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2631__B1 _2429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2891_ _4313_/Q input49/X _2904_/S vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__mux2_8
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2702__B _4122_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3086__A _3099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3512_ _4142_/Q _3308_/A _2767_/A _3490_/A _3504_/X vssd1 vssd1 vccd1 vccd1 _4142_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3443_ _3443_/A vssd1 vssd1 vccd1 vccd1 _4112_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3236__D _3245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4106__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2698__A0 _3291_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2147__C1 _2064_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3814__A _3814_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3374_ _3383_/A _3389_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3375_/A sky130_fd_sc_hd__or3_1
XANTENNA__2162__A2 _2001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2325_ _2301_/X _2302_/X _2324_/X _2304_/X _4361_/Q vssd1 vssd1 vccd1 vccd1 _2325_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4256__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2256_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4067__D _4067_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2187_ _2187_/A _2187_/B vssd1 vssd1 vccd1 vccd1 _2211_/B sky130_fd_sc_hd__nor2_2
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3708__B _4239_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2925__A1 input55/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3724__A _3767_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2689__A0 _3893_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2050__D _2050_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2059__B _2059_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3102__A1 _4202_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3618__B _3635_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4129__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2916__A1 _4107_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2949__S _2949_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output263_A _2738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3634__A _3634_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4279__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3341__A1 _4070_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2144__A2 _2143_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2110_ _2384_/A _2382_/A _2383_/A _2109_/Y vssd1 vssd1 vccd1 vccd1 _2226_/A sky130_fd_sc_hd__o31a_4
X_3090_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3090_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2684__S _3161_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2041_ _2036_/Y _1962_/A _2040_/Y vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__o21ai_2
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3992_ _3992_/A vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2943_ _2943_/A _3447_/B _3442_/C vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__and3_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3809__A _3881_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2713__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2874_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2080__A1 _2204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3247__C _3247_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4350__D _4350_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3544__A _3544_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3426_ _3431_/A _3437_/B _3426_/C vssd1 vssd1 vccd1 vccd1 _3427_/A sky130_fd_sc_hd__or3_1
XFILLER_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3357_ _3369_/A vssd1 vssd1 vccd1 vccd1 _3365_/B sky130_fd_sc_hd__clkbuf_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2308_ _2514_/A vssd1 vssd1 vccd1 vccd1 _2308_/X sky130_fd_sc_hd__buf_4
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3288_ _3320_/A _3288_/B _3323_/C _3317_/C vssd1 vssd1 vccd1 vccd1 _3289_/A sky130_fd_sc_hd__or4_1
X_2239_ _3578_/A _2236_/X _2238_/X vssd1 vssd1 vccd1 vccd1 _2239_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2623__A _2638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2071__B2 _2136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4260__D _4260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2359__C1 _2358_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2374__A2 _2329_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3454__A _3454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input22_A cpu_adr_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3620__C _3624_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3629__A _3629_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2533__A _2533_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2062__A1 _1952_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3067__C _3598_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4170__D _4170_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2590_ _2590_/A _2590_/B _2590_/C _2590_/D vssd1 vssd1 vccd1 vccd1 _2590_/Y sky130_fd_sc_hd__nand4_2
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3364__A _3461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4260_ _4262_/CLK _4260_/D vssd1 vssd1 vccd1 vccd1 _4260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4191_ _4199_/CLK _4191_/D vssd1 vssd1 vccd1 vccd1 _4191_/Q sky130_fd_sc_hd__dfxtp_1
X_3211_ _3211_/A vssd1 vssd1 vccd1 vccd1 _4020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3142_ _3151_/A _3142_/B _3648_/A vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__and3_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2522__C1 _2454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2708__A _2708_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3210_/B _4194_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3602_/C sky130_fd_sc_hd__mux2_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _2024_/A _2072_/B _2081_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__2825__A0 _4302_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4345__D _4345_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2146__C _2210_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3539__A _3546_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3975_ _4369_/Q _3965_/X _2468_/Y _3966_/Y vssd1 vssd1 vccd1 vccd1 _4369_/D sky130_fd_sc_hd__a211o_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3786__D1 _2398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2926_ _3869_/A _4039_/Q _2936_/S vssd1 vssd1 vccd1 vccd1 _3260_/C sky130_fd_sc_hd__mux2_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2857_ _3841_/A _4027_/Q _2905_/S vssd1 vssd1 vccd1 vccd1 _3227_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4080__D _4080_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2447__B1_N _4157_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2788_ _2788_/A vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3553__A1 _3553_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3274__A _3274_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3409_ _3433_/A vssd1 vssd1 vccd1 vccd1 _3429_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4389_ _4389_/CLK _4389_/D vssd1 vssd1 vccd1 vccd1 _4389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3721__B _4247_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3069__A0 _3208_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2337__B _2520_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2277__D1 _2276_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2816__A0 _3823_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4255__D _4255_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3449__A _3457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2029__D1 _2136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2353__A _4152_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2595__A2 _2428_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2072__B _2072_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2503__D _2503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3184__A _3192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output226_A _3133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2528__A _3428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3631__B _3635_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4317__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2962__S _3150_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4165__D _4165_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3359__A _3359_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3760_ _3752_/X _3747_/X _3748_/X _2493_/Y _3757_/X vssd1 vssd1 vccd1 vccd1 _4265_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__2263__A _2346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2035__A1 _2032_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _2715_/A _4126_/Q vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__and2_1
XANTENNA__2586__A2 _2501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__A1 _3769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _4232_/Q _3351_/X _4394_/A _3678_/X _3683_/X vssd1 vssd1 vccd1 vccd1 _4232_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2642_ _2328_/A _2329_/A _4002_/A _2246_/X vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__o211a_1
Xoutput304 _2944_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput315 _2960_/X vssd1 vssd1 vccd1 vccd1 spi_sel_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__3094__A _3094_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2338__A2 _2539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2573_ _2363_/X _2449_/X _2517_/X _2450_/X _4380_/Q vssd1 vssd1 vccd1 vccd1 _2573_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4312_ _4391_/CLK _4312_/D vssd1 vssd1 vccd1 vccd1 _4312_/Q sky130_fd_sc_hd__dfxtp_1
X_4243_ _4264_/CLK _4243_/D vssd1 vssd1 vccd1 vccd1 _4243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3822__A _3822_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4174_ _4177_/CLK _4174_/D vssd1 vssd1 vccd1 vccd1 _4174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3125_ _3135_/A _3125_/B _3635_/C vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__and3_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3541__B _3541_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2510__A2 _2505_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _3192_/C _4189_/Q _3076_/S vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3260__C _3260_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4075__D _4075_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2007_ _2007_/A vssd1 vssd1 vccd1 vccd1 _2160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3471__B1 _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3269__A _3273_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2026__A1 _2204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2577__A2 _2452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _4360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2909_ _4316_/Q input52/X _2940_/S vssd1 vssd1 vccd1 vccd1 _3863_/C sky130_fd_sc_hd__mux2_2
X_3889_ _3889_/A _3893_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__and3_1
XANTENNA__2901__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3526__A1 _3526_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__D1 _3938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3732__A _3748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2348__A _2474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3451__B _3459_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input124_A spi_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A2 _2357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2083__A _2083_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3179__A _3179_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2017__A1 _1962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2568__A2 _2302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3907__A _3907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2530__B _2644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3626__B _3635_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output176_A _2963_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_0_CLK CLK vssd1 vssd1 vccd1 vccd1 clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__3922__D1 _3331_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2957__S _2957_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2258__A _2474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3361__B _3381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2692__S _2949_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3089__A _3099_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3812_ _3884_/A vssd1 vssd1 vccd1 vccd1 _3831_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2008__A1 _2120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3756__A1 _4262_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2559__A2 _2375_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3756__B2 _2466_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3743_ _3727_/X _3729_/X _3732_/X _2338_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _4255_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3239__D _3260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3817__A _3817_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2721__A _2721_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3674_ _3674_/A vssd1 vssd1 vccd1 vccd1 _4224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2440__B _3677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2625_ _2474_/X _2256_/X _2453_/A _2454_/A _2624_/Y vssd1 vssd1 vccd1 vccd1 _2625_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput167 _2642_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput156 _2564_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[20] sky130_fd_sc_hd__buf_2
X_2556_ _4271_/Q vssd1 vssd1 vccd1 vccd1 _2556_/Y sky130_fd_sc_hd__inv_2
Xoutput145 _2460_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput178 _2994_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[11] sky130_fd_sc_hd__buf_2
Xoutput189 _3016_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[21] sky130_fd_sc_hd__buf_2
XANTENNA__3552__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2487_ _2507_/A _3677_/A _2507_/C _2487_/D vssd1 vssd1 vccd1 vccd1 _2487_/Y sky130_fd_sc_hd__nand4_1
XFILLER_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4226_ _4262_/CLK _4226_/D vssd1 vssd1 vccd1 vccd1 _4226_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2495__A1 _2386_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4157_ _4177_/CLK _4157_/D vssd1 vssd1 vccd1 vccd1 _4157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3271__B _3271_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2168__A _2168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3108_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3125_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4088_ _4251_/CLK _4088_/D vssd1 vssd1 vccd1 vccd1 _4088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3039_ _3184_/C _4185_/Q _3157_/S vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3995__A1 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2053__D _2072_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4012__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3727__A _3769_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4162__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__D1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2183__B1 _4345_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3462__A _3586_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2806__A _2828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2238__A1 _2367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__A1 _3952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__B1 _4052_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output293_A _2889_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput25 cpu_adr_i[30] vssd1 vssd1 vccd1 vccd1 _2053_/C sky130_fd_sc_hd__buf_2
XANTENNA__3637__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput14 cpu_adr_i[20] vssd1 vssd1 vccd1 vccd1 _2043_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput36 cpu_dat_i[10] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
Xinput58 cpu_dat_i[30] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
Xinput47 cpu_dat_i[20] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput69 cpu_sel_i[2] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
X_2410_ _4259_/Q vssd1 vssd1 vccd1 vccd1 _2410_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _3390_/A vssd1 vssd1 vccd1 vccd1 _4090_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2174__B1 _2173_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2341_ _2328_/X _2329_/X _3960_/A _2125_/X vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__o211a_2
XANTENNA__3910__A1 _4335_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2687__S _2953_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2272_ _2272_/A _2272_/B input73/X vssd1 vssd1 vccd1 vccd1 _2336_/A sky130_fd_sc_hd__nor3b_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3372__A _3372_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4011_ _4051_/CLK _4011_/D vssd1 vssd1 vccd1 vccd1 _4011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2477__A1 _2475_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2716__A _2716_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2229__A1 _4180_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4035__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4353__D _4353_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1988__B1 _4334_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ input3/X vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__clkinv_2
X_3726_ _2099_/Y _3167_/B _3678_/X _3470_/A vssd1 vssd1 vccd1 vccd1 _4250_/D sky130_fd_sc_hd__a211oi_1
XANTENNA__3547__A _3547_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4185__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2952__A2 _2133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3657_ _3657_/A _3657_/B _3657_/C vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__and3_1
X_2608_ _2638_/A _2638_/B _2638_/C _2608_/D vssd1 vssd1 vccd1 vccd1 _2608_/Y sky130_fd_sc_hd__nand4_2
X_3588_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3609_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2165__B1 _2164_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2539_ _2539_/A vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3901__A1 _3900_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3282__A _3295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__B2 _2398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2468__A1 _2380_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4209_ _4275_/CLK _4209_/D vssd1 vssd1 vccd1 vccd1 _4209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2048__D _2081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2625__D1 _2624_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4263__D _4263_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2640__A1 _2258_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3457__A _3457_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input52_A cpu_dat_i[25] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2156__B1 _3942_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3192__A _3192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2459__A1 _3539_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4058__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3131__S _3144_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output306_A _2788_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3959__A1 _3952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4173__D _4173_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2890_ _2919_/A vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2631__B2 _2430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2631__A1 _2481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2970__S _3335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2271__A _2335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3367__A _3367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3086__B _3089_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3511_ _3511_/A vssd1 vssd1 vccd1 vccd1 _4141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3442_ _3457_/A _3462_/B _3442_/C vssd1 vssd1 vccd1 vccd1 _3443_/A sky130_fd_sc_hd__or3_1
XANTENNA__2698__A1 _4121_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3373_ _3373_/A vssd1 vssd1 vccd1 vccd1 _4083_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2147__B1 _2060_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2429_/A vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__buf_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2255_ _2418_/A vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__buf_4
XFILLER_66_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4348__D _4348_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3830__A _3830_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2186_ _3326_/B _2186_/B _2186_/C _2186_/D vssd1 vssd1 vccd1 vccd1 _2187_/B sky130_fd_sc_hd__nand4b_1
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2446__A _2446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_2_2_0_CLK clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 _4201_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4083__D _4083_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2880__S _2904_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3277__A _3277_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3708__C _3721_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3709_ _3709_/A vssd1 vssd1 vccd1 vccd1 _4239_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3724__B _4249_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2138__B1 _4043_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2689__A1 _4049_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4200__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4258__D _4258_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3740__A _3774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2059__C _2059_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2310__B1 _2309_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2356__A _2356_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4350__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2613__A1 _2319_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2790__S _2826_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2091__A _3489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3187__A _3187_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3618__C _3618_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3915__A _3915_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output256_A _2725_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3341__A2 _3331_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4168__D _4168_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3650__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2040_ _4347_/Q _2012_/B _2038_/Y _2152_/A vssd1 vssd1 vccd1 vccd1 _2040_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ _3991_/A vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2942_ _3267_/B _4112_/Q _2942_/S vssd1 vssd1 vccd1 vccd1 _3442_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2604__A1 _2423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2713__B _4127_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2873_ _2873_/A vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3097__A _3097_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2080__A2 _2018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3247__D _3260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3825__A _3897_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4223__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3425_ _3425_/A vssd1 vssd1 vccd1 vccd1 _4105_/D sky130_fd_sc_hd__clkbuf_1
X_3356_ _3591_/A vssd1 vssd1 vccd1 vccd1 _3470_/A sky130_fd_sc_hd__buf_4
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__D _4078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2307_ _2224_/X _2245_/X _2306_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__o211a_2
XANTENNA__2875__S _2885_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3287_ _3287_/A vssd1 vssd1 vccd1 vccd1 _4049_/D sky130_fd_sc_hd__clkbuf_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__A _3562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2238_ _2367_/A _2335_/A _4283_/Q vssd1 vssd1 vccd1 vccd1 _2238_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4373__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2047__B1_N _4345_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2169_ _2167_/Y _3902_/A _2013_/Y _2153_/C vssd1 vssd1 vccd1 vccd1 _2169_/Y sky130_fd_sc_hd__o211ai_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2623__B _2638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2359__B1 _2246_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3735__A _3771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2785__S _3790_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3470__A _3470_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input15_A cpu_adr_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2814__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3629__B _3633_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2062__A2 _2007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4246__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3645__A _3645_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2770__A0 _4293_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4190_ _4286_/CLK _4190_/D vssd1 vssd1 vccd1 vccd1 _4190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3210_ _3224_/A _3210_/B _3224_/C _3219_/D vssd1 vssd1 vccd1 vccd1 _3211_/A sky130_fd_sc_hd__or4_1
X_3141_ _3260_/C _4213_/Q _3147_/S vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2522__B1 _2453_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3380__A _3444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3089_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_95_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2023_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__buf_4
XANTENNA__2825__A1 input37/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2724__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3974_ _3974_/A vssd1 vssd1 vccd1 vccd1 _4368_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3539__B _3539_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3786__C1 _3938_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2925_ _4319_/Q input55/X _2935_/S vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__mux2_4
XANTENNA__4361__D _4361_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2856_ _2958_/S vssd1 vssd1 vccd1 vccd1 _2905_/S sky130_fd_sc_hd__buf_2
XANTENNA__3538__C1 _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2787_ _2799_/A _2812_/B _3376_/A vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__and3_2
XANTENNA__3553__A2 _3365_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3408_ _3408_/A vssd1 vssd1 vccd1 vccd1 _4098_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3710__C1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4388_ _4388_/CLK _4388_/D vssd1 vssd1 vccd1 vccd1 _4388_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input7_A cpu_adr_i[14] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3339_ _3339_/A vssd1 vssd1 vccd1 vccd1 _4069_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3290__A _3707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3721__C _3721_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3069__A1 _4193_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2277__C1 _2409_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4119__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2816__A1 _4020_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2337__C _2520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2029__C1 _2015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3449__B _3462_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4269__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3777__C1 _3774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4271__D _4271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3529__C1 _3562_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2072__C _2078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3465__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3184__B _3199_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3701__C1 _3683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3631__C _3631_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output219_A _3111_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3768__C1 _3755_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2035__A2 _1962_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2710_ _2710_/A vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3783__A2 _3764_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4181__D _4181_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _3690_/A vssd1 vssd1 vccd1 vccd1 _4231_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2436__B_N _2383_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3375__A _3375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2641_ _3562_/B _2526_/A _2636_/Y _2640_/Y vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__o211ai_4
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput305 _2781_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput316 _4395_/X vssd1 vssd1 vccd1 vccd1 spi_stb_o sky130_fd_sc_hd__buf_2
X_2572_ _2572_/A1 _2444_/X _2514_/X _2445_/X _2571_/Y vssd1 vssd1 vccd1 vccd1 _3554_/B
+ sky130_fd_sc_hd__a41oi_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4311_ _4371_/CLK _4311_/D vssd1 vssd1 vccd1 vccd1 _4311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4242_ _4264_/CLK _4242_/D vssd1 vssd1 vccd1 vccd1 _4242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2719__A _2719_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4173_ _4180_/CLK _4173_/D vssd1 vssd1 vccd1 vccd1 _4173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3124_ _3245_/B _4208_/Q _3144_/S vssd1 vssd1 vccd1 vccd1 _3635_/C sky130_fd_sc_hd__mux2_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3055_ _3657_/B vssd1 vssd1 vccd1 vccd1 _3070_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3260__D _3260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4356__D _4356_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2006_ input9/X vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3471__B2 _3469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3471__A1 _4122_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2454__A _2454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3759__C1 _3755_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3957_ _3957_/A _3973_/B _3963_/C vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__and3_1
XANTENNA__3269__B _3279_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2026__A2 _2018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2908_ _2908_/A vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2431__C1 _4366_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4091__D _4091_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2982__B1 _3673_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _3888_/A vssd1 vssd1 vccd1 vccd1 _4326_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2901__B _2901_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2839_ _3834_/C _4024_/Q _2886_/S vssd1 vssd1 vccd1 vccd1 _3219_/B sky130_fd_sc_hd__mux2_4
XANTENNA__3285__A _3692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3526__A2 _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__C1 _3909_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3451__C _3455_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4266__D _4266_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input117_A spi_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4091__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2083__B _2083_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2017__A2 _2012_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input82_A gpio_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3195__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2530__C _2530_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3626__C _3626_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3922__C1 _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output169_A _2327_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3642__B _3659_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3150__A0 _3267_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2539__A _2539_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__S _3147_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3361__C _3376_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4176__D _4176_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2274__A _2638_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3089__B _3089_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3811_ _3811_/A vssd1 vssd1 vccd1 vccd1 _4294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2008__A2 _2160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3756__A2 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3742_ _4254_/Q _3734_/X _3735_/X input99/X _3738_/X vssd1 vssd1 vccd1 vccd1 _4254_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3673_ _3798_/A _3673_/B _3673_/C vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__or3_1
XANTENNA__3817__B _3821_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2624_ _2622_/Y _2366_/A _2623_/Y vssd1 vssd1 vccd1 vccd1 _2624_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__2440__C _2507_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3913__C1 _3912_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2177__D1 _2136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput168 _2649_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput157 _2570_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[21] sky130_fd_sc_hd__buf_2
X_2555_ _2512_/X _2513_/X _2554_/Y _2524_/X vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3833__A _3881_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput146 _2470_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput179 _2996_/X vssd1 vssd1 vccd1 vccd1 gpio_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2486_ _4264_/Q vssd1 vssd1 vccd1 vccd1 _2486_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3552__B _3552_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2449__A _2474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3141__A0 _3260_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4225_ _4225_/CLK _4225_/D vssd1 vssd1 vccd1 vccd1 _4225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _4172_/CLK _4156_/D vssd1 vssd1 vccd1 vccd1 _4156_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3271__C _3276_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3107_ _3107_/A vssd1 vssd1 vccd1 vccd1 _3107_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2495__A2 _2424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4086__D _4086_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4225_/CLK _4087_/D vssd1 vssd1 vccd1 vccd1 _4087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3038_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3044_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3995__A2 _3992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2184__A _2184_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2912__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2955__A0 _3178_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4307__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__C1 _3938_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2183__A1 _2121_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3462__B _3462_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2078__B _2078_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2806__B _2812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2238__A2 _2335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__A2 _3955_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__A1 _1993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3918__A _3918_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2946__A0 _3792_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 cpu_adr_i[31] vssd1 vssd1 vccd1 vccd1 _2061_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output286_A _2853_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput15 cpu_adr_i[21] vssd1 vssd1 vccd1 vccd1 _2182_/A sky130_fd_sc_hd__buf_2
Xinput37 cpu_dat_i[11] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput59 cpu_dat_i[31] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_4
Xinput48 cpu_dat_i[21] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2968__S _3150_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3653__A _3653_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2174__A1 _2171_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _3530_/B _2255_/X _2333_/Y _2339_/Y vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__o211ai_4
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3910__A2 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2271_ _2335_/A vssd1 vssd1 vccd1 vccd1 _2590_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__2269__A _2344_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3372__B _3381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4010_ _4051_/CLK _4010_/D vssd1 vssd1 vccd1 vccd1 _4010_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2477__A2 _2366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2229__A2 _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1988__A1 _1930_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3828__A _3876_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2732__A _2732_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2937__A0 _3265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _4335_/Q _2182_/B _1983_/Y _2137_/A _1985_/X vssd1 vssd1 vccd1 vccd1 _1986_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3725_ _3725_/A vssd1 vssd1 vccd1 vccd1 _4249_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3039__S _3157_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3656_ _3656_/A vssd1 vssd1 vccd1 vccd1 _4216_/D sky130_fd_sc_hd__clkbuf_1
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _4188_/D sky130_fd_sc_hd__clkbuf_1
X_2607_ _4277_/Q vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2165__A1 _2028_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2538_ _4269_/Q vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3901__A2 _1998_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4208_ _4280_/CLK _4208_/D vssd1 vssd1 vccd1 vccd1 _4208_/Q sky130_fd_sc_hd__dfxtp_1
X_2469_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__A2 _2464_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4139_ _4141_/CLK _4139_/D vssd1 vssd1 vccd1 vccd1 _4139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4394__A _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2907__A _2917_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2625__C1 _2454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3738__A _3772_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2640__A2 _2256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3457__B _3462_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3473__A _3516_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2156__B2 _2136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2089__A _2529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A cpu_dat_i[19] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3192__B _3199_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3105__A0 _3234_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2459__A2 _2362_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output201_A _2971_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2616__C1 _4385_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3959__A2 _3955_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2631__A2 _2501_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2552__A _2552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3648__A _3648_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3367__B _3381_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3510_ _3510_/A _4141_/Q _3657_/C vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__and3_1
XANTENNA__3086__C _3609_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3462_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3383__A _3383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2698__S _2947_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2147__A1 _3346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3372_ _3372_/A _3381_/B _3376_/C vssd1 vssd1 vccd1 vccd1 _3373_/A sky130_fd_sc_hd__and3_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2323_ _4254_/Q _2322_/X _2298_/X input99/X vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_69_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2254_ _2254_/A1 _2090_/A _2248_/X _2421_/A _2253_/Y vssd1 vssd1 vccd1 vccd1 _3522_/B
+ sky130_fd_sc_hd__a41oi_4
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2727__A _2727_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2185_ _4065_/Q _1977_/X _2184_/Y vssd1 vssd1 vccd1 vccd1 _2186_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4364__D _4364_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4152__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3558__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3708__D _3711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1969_ _2093_/A vssd1 vssd1 vccd1 vccd1 _3332_/A sky130_fd_sc_hd__clkbuf_2
X_3708_ _3717_/A _4239_/Q _3721_/C _3711_/D vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__and4_1
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3639_ _3639_/A vssd1 vssd1 vccd1 vccd1 _4209_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3724__C _3724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3293__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2138__A1 _2136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2637__A _4281_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2310__A1 _2310_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4274__D _4274_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2356__B _2356_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2613__A2 _2248_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3468__A _3468_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2372__A _2579_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4025__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output249_A _2710_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output151_A _2525_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3650__B _3659_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4175__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4184__D _4184_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2981__S _3150_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3990_/A vssd1 vssd1 vccd1 vccd1 _4380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2604__A2 _2446_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2941_ _3877_/C _4042_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _3267_/B sky130_fd_sc_hd__mux2_4
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2282__A _2543_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3378__A _3383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2872_ _2888_/A _2872_/B _3410_/A vssd1 vssd1 vccd1 vccd1 _2873_/A sky130_fd_sc_hd__and3_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4002__A _4002_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3424_ _3424_/A _3429_/B _3424_/C vssd1 vssd1 vccd1 vccd1 _3425_/A sky130_fd_sc_hd__and3_1
XANTENNA__4359__D _4359_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3355_ _3355_/A vssd1 vssd1 vccd1 vccd1 _4077_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3841__A _3841_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2306_ _2281_/X _2291_/Y _2293_/X _2299_/Y _2305_/Y vssd1 vssd1 vccd1 vccd1 _2306_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_58_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3286_ _3328_/B _3689_/D _3286_/C _3286_/D vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__and4_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__B _3560_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ _2237_/A vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__clkbuf_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4094__D _4094_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2168_/A vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__buf_2
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2099_ _4250_/Q vssd1 vssd1 vccd1 vccd1 _2099_/Y sky130_fd_sc_hd__inv_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2891__S _2904_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2056__B1 _2134_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2192__A _2782_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3288__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2623__C _2638_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2359__A1 _2328_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4048__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4269__D _4269_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4198__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2367__A _2367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2598__A1 _2319_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3198__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3629__C _3648_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output199_A _3035_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2830__A _3489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3926__A _3926_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_CLK clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2107__B1_N _4285_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2770__A1 input57/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4179__D _4179_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3140_ _3140_/A vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2522__A1 _2474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3661__A _3661_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3071_ _3071_/A vssd1 vssd1 vccd1 vccd1 _3071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2022_ _2022_/A vssd1 vssd1 vccd1 vccd1 _2081_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2724__B _4132_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3786__B1 _2238_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3973_ _3973_/A _3973_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__and3_1
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2924_ _2924_/A vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2855_ _4307_/Q input42/X _2904_/S vssd1 vssd1 vccd1 vccd1 _3841_/A sky130_fd_sc_hd__mux2_8
XANTENNA__2740__A _2748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3538__B1 _2437_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3836__A _3884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2786_ _3192_/C _4085_/Q _2955_/S vssd1 vssd1 vccd1 vccd1 _3376_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3553__A3 _3544_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4340__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3407_ _3407_/A _3413_/B _3407_/C vssd1 vssd1 vccd1 vccd1 _3408_/A sky130_fd_sc_hd__or3_1
X_4387_ _4389_/CLK _4387_/D vssd1 vssd1 vccd1 vccd1 _4387_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2886__S _2886_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4089__D _4089_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3710__B1 _3696_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3571__A _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3338_ _2158_/A _3488_/A _3724_/D _3724_/C vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__and4b_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3721__D _3724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3269_ _3273_/A _3279_/B _3269_/C _3286_/D vssd1 vssd1 vccd1 vccd1 _3270_/A sky130_fd_sc_hd__and4_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2187__A _2187_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2277__B1 _2408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2337__D _2337_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2029__B1 _2028_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3449__C _3449_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3777__B1 _2591_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3529__B1 _2320_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2072__D _2078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2650__A _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3184__C _3184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3481__A _3481_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3701__B1 _3696_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2504__A1 _2287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4213__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3768__B1 _3754_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3783__A3 _3748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3656__A _3656_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2640_ _2258_/X _2256_/X _2453_/A _2454_/A _2639_/Y vssd1 vssd1 vccd1 vccd1 _2640_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4363__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput306 _2788_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput317 _2194_/X vssd1 vssd1 vccd1 vccd1 spi_we_o sky130_fd_sc_hd__buf_2
X_2571_ _2423_/A _2446_/X _4169_/Q vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__a21boi_1
X_4310_ _4371_/CLK _4310_/D vssd1 vssd1 vccd1 vccd1 _4310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4241_ _4264_/CLK _4241_/D vssd1 vssd1 vccd1 vccd1 _4241_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3391__A _3391_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4172_ _4172_/CLK _4172_/D vssd1 vssd1 vccd1 vccd1 _4172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _3123_/A vssd1 vssd1 vccd1 vccd1 _3123_/X sky130_fd_sc_hd__clkbuf_1
X_3054_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__buf_2
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__A _2737_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2005_ _2146_/B _3303_/B _2005_/C _2098_/B vssd1 vssd1 vccd1 vccd1 _2129_/A sky130_fd_sc_hd__nand4b_4
XANTENNA__3471__A2 _3350_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4372__D _4372_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3759__B1 _3754_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3956_ _3952_/X _3955_/X _2306_/Y vssd1 vssd1 vccd1 vccd1 _4359_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__3269__C _3269_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2907_ _2917_/A _2928_/B _3424_/A vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__and3_1
XANTENNA__2431__B1 _2429_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2982__A1 _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3566__A _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _3895_/A _3935_/B _3887_/C vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__or3_1
XANTENNA__2901__C _3422_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2838_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2886_/S sky130_fd_sc_hd__buf_2
X_2769_ _3489_/A vssd1 vssd1 vccd1 vccd1 _2799_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3526__A3 _3524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__B1 _2078_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2498__B1 _2497_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4236__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2670__A0 _3887_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4282__D _4282_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4386__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2083__C _2083_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2017__A3 _2013_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2380__A _2380_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3195__B _3195_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_27_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4326_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input75_A gpio_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3922__B1 _2013_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__C _3642_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2489__B1 _2488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3150__A1 _4216_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output231_A _3050_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3150__S _3150_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2661__A0 _4325_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3089__C _3611_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4192__D _4192_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3823_/A _3829_/B _3810_/C vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__or3_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3741_ _3727_/X _3729_/X _3732_/X _2315_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _4253_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3386__A _3386_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3672_ _3672_/A vssd1 vssd1 vccd1 vccd1 _4223_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_18_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4275_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3817__C _3831_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2623_ _2638_/A _2638_/B _2638_/C _2623_/D vssd1 vssd1 vccd1 vccd1 _2623_/Y sky130_fd_sc_hd__nand4_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2440__D _2440_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2554_ _2281_/X _2550_/Y _2293_/X _2551_/Y _2553_/Y vssd1 vssd1 vccd1 vccd1 _2554_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4109__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3913__B1 _3911_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2177__C1 _1973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput158 _2580_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput147 _2480_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2485_ _2283_/X _2483_/X _2484_/Y vssd1 vssd1 vccd1 vccd1 _2485_/Y sky130_fd_sc_hd__a21oi_2
Xoutput169 _2327_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[3] sky130_fd_sc_hd__buf_2
X_4224_ _4262_/CLK _4224_/D vssd1 vssd1 vccd1 vccd1 _4224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4259__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4155_ _4389_/CLK _4155_/D vssd1 vssd1 vccd1 vccd1 _4155_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3141__A1 _4213_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4367__D _4367_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3271__D _3271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3106_ _3117_/A _3106_/B _3624_/A vssd1 vssd1 vccd1 vccd1 _3107_/A sky130_fd_sc_hd__and3_1
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4086_ _4251_/CLK _4086_/D vssd1 vssd1 vccd1 vccd1 _4086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2465__A _4262_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2184__B _2184_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2652__A0 _4324_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2912__B _2928_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2955__A1 _4079_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3939_ _2061_/Y _3902_/A _2062_/Y vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3904__B1 _2002_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2183__A2 _2160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3462__C _3462_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4277__D _4277_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2340__C1 _2339_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2078__C _2078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2891__A0 _4313_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2806__C _3383_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2375__A _2375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__A2 _1996_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3918__B _3942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 cpu_adr_i[22] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
XANTENNA__2946__A1 _4007_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 cpu_adr_i[3] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output181_A _3000_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput49 cpu_dat_i[22] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 cpu_dat_i[12] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output279_A _4395_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3653__B _3661_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2174__A2 _2153_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2270_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3372__C _3376_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4187__D _4187_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_7_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4172_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2882__A0 _3239_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2285__A _2531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2095__D1 _3301_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1988__A2 _2141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1985_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__clkbuf_4
X_3724_ _3767_/A _4249_/Q _3724_/C _3724_/D vssd1 vssd1 vccd1 vccd1 _3725_/A sky130_fd_sc_hd__and4_1
XANTENNA__2937__A1 _4111_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3655_ _3659_/A _3659_/B _3655_/C vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__or3_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2606_ _2427_/A _2449_/X _2517_/X _2450_/X _4384_/Q vssd1 vssd1 vccd1 vccd1 _2606_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3844__A _3844_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3586_ _3586_/A _3586_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__or3_1
XANTENNA__4081__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2165__A2 _2001_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2537_ _2512_/X _2513_/X _2246_/X _2536_/Y vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__o211a_1
X_2468_ _2380_/X _2464_/Y _2467_/X _2398_/X vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__2570__C1 _2524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4207_ _4275_/CLK _4207_/D vssd1 vssd1 vccd1 vccd1 _4207_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4097__D _4097_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2399_ _2380_/X _2389_/Y _2397_/X _2398_/X vssd1 vssd1 vccd1 vccd1 _2399_/Y sky130_fd_sc_hd__o22ai_4
X_4138_ _4141_/CLK _4138_/D vssd1 vssd1 vccd1 vccd1 _4138_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2907__B _2928_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2195__A _4250_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4069_ _4380_/CLK _4069_/D vssd1 vssd1 vccd1 vccd1 _4069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2625__B1 _2453_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2923__A _2943_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3457__C _3457_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3754__A _3771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3192__C _3192_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3105__A1 _4203_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input38_A cpu_dat_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2616__B1 _2324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3648__B _3661_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3367__C _3376_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2979__S _3157_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3664__A _3798_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _3440_/A vssd1 vssd1 vccd1 vccd1 _4111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3371_ _3371_/A vssd1 vssd1 vccd1 vccd1 _4082_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3383__B _3389_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2147__A2 _3346_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2322_ _3720_/A vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__buf_6
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2253_ _2644_/A _2424_/A _4147_/Q vssd1 vssd1 vccd1 vccd1 _2253_/Y sky130_fd_sc_hd__a21boi_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2855__A0 _4307_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2184_ _2184_/A _2184_/B _2184_/C vssd1 vssd1 vccd1 vccd1 _2184_/Y sky130_fd_sc_hd__nand3_1
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3839__A _3847_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2743__A _2743_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3558__B _3558_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4380__D _4380_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1968_ _4056_/Q vssd1 vssd1 vccd1 vccd1 _1968_/Y sky130_fd_sc_hd__inv_2
X_3707_ _3707_/A vssd1 vssd1 vccd1 vccd1 _3721_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3574__A _3574_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3638_ _3638_/A _3661_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__and3_1
XANTENNA__3724__D _3724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3569_ _3569_/A _3584_/B _3657_/A vssd1 vssd1 vccd1 vccd1 _3570_/A sky130_fd_sc_hd__and3_1
XANTENNA__3293__B _3335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2138__A2 _3942_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2918__A _2918_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2846__A0 _3221_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2310__A2 _2090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2356__C _2356_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2653__A _2662_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4290__D _4290_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2828__A _2828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output144_A _2279_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3650__C _3650_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2837__A0 _4304_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output311_A _2819_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3659__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _4322_/Q input59/X _2940_/S vssd1 vssd1 vccd1 vccd1 _3877_/C sky130_fd_sc_hd__mux2_1
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3378__B _3389_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2871_ _3234_/C _4099_/Q _2916_/S vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__mux2_4
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3394__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3423_ _3423_/A vssd1 vssd1 vccd1 vccd1 _4104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4002__B _4002_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2525__C1 _2524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3354_ _3354_/A _3774_/A _3376_/C vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__and3_1
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2738__A _2738_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2305_ _2301_/X _2302_/X _2303_/X _2304_/X _4359_/Q vssd1 vssd1 vccd1 vccd1 _2305_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3285_ _3692_/A vssd1 vssd1 vccd1 vccd1 _3689_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__3841__B _3845_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2236_ _2964_/A _2139_/Y _2213_/Y vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__o21a_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4375__D _4375_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2167_ _2167_/A vssd1 vssd1 vccd1 vccd1 _2167_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2098_ _2098_/A _2098_/B _2098_/C _2098_/D vssd1 vssd1 vccd1 vccd1 _2112_/B sky130_fd_sc_hd__nand4_4
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3569__A _3569_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2056__A1 _3938_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3288__B _3288_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2623__D _2623_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2359__A2 _2329_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4285__D _4285_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2383__A _2383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2047__A1 _2120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2598__A2 _2248_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4142__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output261_A _2734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3942__A _3942_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3153__S _3157_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2522__A2 _2452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3661__B _3661_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _3081_/A _3070_/B _3600_/A vssd1 vssd1 vccd1 vccd1 _3071_/A sky130_fd_sc_hd__and3_1
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4195__D _4195_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2021_ _2078_/B vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4292__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2293__A _2509_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3389__A _3407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3786__A1 _3734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3972_ _4002_/C vssd1 vssd1 vccd1 vccd1 _3996_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2923_ _2943_/A _2928_/B _3431_/C vssd1 vssd1 vccd1 vccd1 _2924_/A sky130_fd_sc_hd__and3_1
X_2854_ _2957_/S vssd1 vssd1 vccd1 vccd1 _2904_/S sky130_fd_sc_hd__buf_4
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2740__B _4139_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3538__A1 _2436_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2785_ _3813_/A _4015_/Q _3790_/A vssd1 vssd1 vccd1 vccd1 _3192_/C sky130_fd_sc_hd__mux2_4
XANTENNA__3852__A _3876_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4386_ _4388_/CLK _4386_/D vssd1 vssd1 vccd1 vccd1 _4386_/Q sky130_fd_sc_hd__dfxtp_1
X_3406_ _3406_/A vssd1 vssd1 vccd1 vccd1 _4097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3710__A1 _4240_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3710__B2 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3337_ _3800_/A vssd1 vssd1 vccd1 vccd1 _3724_/C sky130_fd_sc_hd__buf_6
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3268_ _3268_/A vssd1 vssd1 vccd1 vccd1 _4042_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2187__B _2187_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2219_ _2257_/A vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__2277__A1 _2262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3199_ _3221_/A _3199_/B _3199_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3200_/A sky130_fd_sc_hd__and4_1
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3299__A _3343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2029__A1 _4341_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3777__A1 _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4015__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3529__A1 _3529_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4165__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__D1 _3938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3184__D _3208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3701__A1 _4236_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3701__B2 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2504__A2 _2424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2378__A _2552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A cpu_adr_i[26] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3002__A _3010_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3768__A1 _4270_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3768__B2 input84/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2841__A _2859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput307 _2793_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[5] sky130_fd_sc_hd__buf_2
X_2570_ _2512_/X _2513_/X _2569_/Y _2524_/X vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3672__A _3672_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4264_/CLK _4240_/D vssd1 vssd1 vccd1 vccd1 _4240_/Q sky130_fd_sc_hd__dfxtp_1
X_4171_ _4177_/CLK _4171_/D vssd1 vssd1 vccd1 vccd1 _4171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2288__A _2446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3391__B _3405_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3135_/A _3125_/B _3633_/A vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__and3_1
XFILLER_95_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3053_ _3053_/A vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4038__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1920__A _1934_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2004_ _3294_/C _3294_/B _2145_/C _2145_/D vssd1 vssd1 vccd1 vccd1 _2098_/B sky130_fd_sc_hd__and4_2
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2735__B _4137_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3759__A1 _4264_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3759__B2 _2487_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3955_ _3992_/A vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3269__D _3286_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2751__A _2751_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4188__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2431__B2 _2430_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2431__A1 _2427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2906_ _3247_/C _4105_/Q _2916_/S vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3847__A _3847_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2982__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3886_ _3886_/A vssd1 vssd1 vccd1 vccd1 _4325_/D sky130_fd_sc_hd__clkbuf_1
X_2837_ _4304_/Q input39/X _2885_/S vssd1 vssd1 vccd1 vccd1 _3834_/C sky130_fd_sc_hd__mux2_2
X_2768_ _2768_/A vssd1 vssd1 vccd1 vccd1 _2768_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2699_ _2677_/X _2680_/X _3466_/A vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2897__S _2940_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__A1 _4349_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3582__A _3586_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2498__A1 _2419_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2198__A _2349_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4369_ _4390_/CLK _4369_/D vssd1 vssd1 vccd1 vccd1 _4369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3998__A1 _3991_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_CLK clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2670__A1 _4046_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3757__A _3774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2083__D _2083_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3195__C _3195_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input68_A cpu_sel_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__A1 _2167_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3492__A _3492_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1933__B1 _4338_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2489__B2 _2398_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2489__A1 _2380_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output224_A _3126_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2836__A _2896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2110__B1 _2109_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2661__A1 input13/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4330__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3740_ _3774_/A vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3667__A _3667_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3386__B _3405_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3671_ _3671_/A _3796_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__and3_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _4279_/Q vssd1 vssd1 vccd1 vccd1 _2622_/Y sky130_fd_sc_hd__inv_2
X_2553_ _2301_/X _2302_/X _2324_/X _2552_/X _4377_/Q vssd1 vssd1 vccd1 vccd1 _2553_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3913__A1 input5/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2177__B1 _2176_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput159 _2588_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput148 _2490_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2484_ _2287_/X _3468_/A _4160_/Q vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4223_ _4286_/CLK _4223_/D vssd1 vssd1 vccd1 vccd1 _4223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4154_ _4172_/CLK _4154_/D vssd1 vssd1 vccd1 vccd1 _4154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2746__A _2748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3105_ _3234_/C _4203_/Q _3112_/S vssd1 vssd1 vccd1 vccd1 _3624_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4085_ _4085_/CLK _4085_/D vssd1 vssd1 vccd1 vccd1 _4085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3036_ _3036_/A _4249_/Q vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__and2_1
XANTENNA__4383__D _4383_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2184__C _2184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2652__A1 input2/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3577__A _3577_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2481__A _3730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2912__C _3426_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3938_ _3938_/A _3938_/B _3938_/C _3938_/D vssd1 vssd1 vccd1 vccd1 _4354_/D sky130_fd_sc_hd__nand4_1
X_3869_ _3869_/A _3869_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__and3_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3904__A1 input33/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4203__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2656__A _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2340__B1 _2333_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2078__D _2078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input122_A spi_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2891__A1 input49/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4353__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4293__D _4293_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3487__A _3487_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2391__A _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3918__C _3940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput17 cpu_adr_i[23] vssd1 vssd1 vccd1 vccd1 _2037_/A sky130_fd_sc_hd__clkbuf_2
Xinput28 cpu_adr_i[4] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
Xinput39 cpu_dat_i[13] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2613__B1_N _4174_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output174_A _2433_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3653__C _3675_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__A _3950_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2882__A1 _4101_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2634__A1 _2423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2095__C1 _1990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3397__A _3397_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1984_ _2055_/B vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__buf_2
X_3723_ _4248_/Q _3167_/B _3044_/A _3697_/A _3470_/A vssd1 vssd1 vccd1 vccd1 _4248_/D
+ sky130_fd_sc_hd__a221o_1
X_3654_ _3654_/A vssd1 vssd1 vccd1 vccd1 _4215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4226__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2605_ _2605_/A1 _2444_/X _2514_/X _2445_/X _2604_/Y vssd1 vssd1 vccd1 vccd1 _3558_/B
+ sky130_fd_sc_hd__a41oi_4
X_3585_ _3585_/A vssd1 vssd1 vccd1 vccd1 _4187_/D sky130_fd_sc_hd__clkbuf_1
X_2536_ _2526_/X _2532_/Y _2509_/X _2534_/Y _2535_/Y vssd1 vssd1 vccd1 vccd1 _2536_/Y
+ sky130_fd_sc_hd__o221ai_4
X_2467_ _2465_/Y _2411_/X _2466_/Y vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__o21a_4
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2570__B1 _2569_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4378__D _4378_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4206_ _4280_/CLK _4206_/D vssd1 vssd1 vccd1 vccd1 _4206_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4376__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3860__A _3884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _2509_/A vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__buf_6
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2156__A2_N _4070_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4137_ _4141_/CLK _4137_/D vssd1 vssd1 vccd1 vccd1 _4137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2907__C _3424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2476__A _2575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4068_ _4391_/CLK _4068_/D vssd1 vssd1 vccd1 vccd1 _4068_/Q sky130_fd_sc_hd__dfxtp_1
X_3019_ _3021_/A _4241_/Q vssd1 vssd1 vccd1 vccd1 _3020_/A sky130_fd_sc_hd__and2_1
XANTENNA__2625__A1 _2474_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2923__B _2928_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3100__A _3100_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2389__B1 _2388_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2561__B1 _2560_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3192__D _3208_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4288__D _4288_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2386__A _2644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3988__B1_N _2569_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2616__A1 _2407_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2616__B2 _2552_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3010__A _3010_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3648__C _3648_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4249__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output291_A _2768_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3945__A _3945_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3664__B _3673_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3370_ _3383_/A _3389_/B _3370_/C vssd1 vssd1 vccd1 vccd1 _3371_/A sky130_fd_sc_hd__or3_1
XANTENNA__3383__C _3383_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2321_ _3529_/A1 _2283_/X _2286_/X _2320_/Y vssd1 vssd1 vccd1 vccd1 _2321_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__4198__D _4198_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3680__A _3680_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2252_ _2514_/A vssd1 vssd1 vccd1 vccd1 _2424_/A sky130_fd_sc_hd__buf_2
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__C1 _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2296__A _2367_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2855__A1 input42/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2183_ _2121_/A _2160_/X _4345_/Q vssd1 vssd1 vccd1 vccd1 _2184_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3839__B _3853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2462__C _2462_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3706_ _4238_/Q _3695_/X _3696_/X _3697_/X _3705_/X vssd1 vssd1 vccd1 vccd1 _4238_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3855__A _3855_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1967_ _2207_/A _2207_/B _3308_/C _1967_/D vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__nand4_1
XANTENNA__2791__A0 _3195_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3574__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3066__S _3073_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3637_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3661_/B sky130_fd_sc_hd__buf_2
XANTENNA__2078__A_N input19/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3568_ _3720_/A vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3293__C _3707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2519_ _4267_/Q vssd1 vssd1 vccd1 vccd1 _2519_/Y sky130_fd_sc_hd__inv_2
X_3499_ _3510_/A _4135_/Q _3502_/C vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__and3_1
XANTENNA__3590__A _3590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2846__A1 _4095_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2310__A3 _2308_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2934__A _2934_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3559__C1 _3547_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3765__A _3765_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2534__B1 _3771_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input50_A cpu_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2828__B _2841_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_19_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2837__A1 input39/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3005__A _3005_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output304_A _2944_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3659__B _3659_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4071__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3378__C _3378_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2470__C1 _2469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2870_ _3197_/A vssd1 vssd1 vccd1 vccd1 _2916_/S sky130_fd_sc_hd__buf_2
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3675__A _3675_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2222__C1 _4390_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3394__B _3413_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3422_ _3431_/A _3437_/B _3422_/C vssd1 vssd1 vccd1 vccd1 _3423_/A sky130_fd_sc_hd__or3_1
XANTENNA__4002__C _4002_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2525__B1 _3982_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3444_/A vssd1 vssd1 vccd1 vccd1 _3376_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1923__A _1923_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2304_/X sky130_fd_sc_hd__buf_2
XFILLER_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3841__C _3855_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3284_ _3284_/A vssd1 vssd1 vccd1 vccd1 _4048_/D sky130_fd_sc_hd__clkbuf_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2235_ _2638_/A _2335_/A vssd1 vssd1 vccd1 vccd1 _3578_/A sky130_fd_sc_hd__nand2_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2166_ _4061_/Q _1977_/X _2165_/Y vssd1 vssd1 vccd1 vccd1 _2175_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2754__A _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2097_ _1949_/Y _2093_/X _1962_/Y _2207_/D vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3789__C1 _3566_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__B _3584_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2056__A2 _3938_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2461__C1 _4369_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4391__D _4391_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3288__C _3323_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2999_ _2999_/A _4232_/Q vssd1 vssd1 vccd1 vccd1 _3000_/A sky130_fd_sc_hd__and2_1
XANTENNA__3585__A _3585_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2764__A0 _3805_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3713__C1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2516__B1 _2515_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2929__A _2929_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4094__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2047__A2 _2141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input98_A gpio_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3495__A _3516_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3942__B _3942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output254_A _2721_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3661__C _3675_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2020_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2024_/A sky130_fd_sc_hd__inv_2
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2574__A _4273_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3389__B _3389_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3971_ _4367_/Q _3965_/X _2442_/Y _3966_/Y vssd1 vssd1 vccd1 vccd1 _4367_/D sky130_fd_sc_hd__a211o_1
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ _3257_/B _4108_/Q _2942_/S vssd1 vssd1 vccd1 vccd1 _3431_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3786__A2 _2236_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2443__C1 _2373_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2853_ _2853_/A vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3538__A2 _3536_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2784_ _4295_/Q input61/X _3907_/A vssd1 vssd1 vccd1 vccd1 _3813_/A sky130_fd_sc_hd__mux2_4
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2749__A _2749_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4385_ _4389_/CLK _4385_/D vssd1 vssd1 vccd1 vccd1 _4385_/Q sky130_fd_sc_hd__dfxtp_1
X_3405_ _3405_/A _3405_/B _3424_/C vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__and3_1
XANTENNA__3710__A2 _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3336_ input1/X vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__buf_4
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__D _4386_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3276_/A _3267_/B _3276_/C _3271_/D vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__or4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2218_ _2346_/A vssd1 vssd1 vccd1 vccd1 _2452_/A sky130_fd_sc_hd__buf_2
XANTENNA__2277__A2 _2375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3221_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2149_ _2662_/A _2148_/Y _2083_/A vssd1 vssd1 vccd1 vccd1 _2158_/A sky130_fd_sc_hd__o21a_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3299__B _3326_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2029__A2 _1970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3777__A2 _3764_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3529__A2 _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3934__C1 _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2659__A _2659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3701__A2 _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__D1 _2369_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4296__D _4296_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2394__A _2638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input13_A cpu_adr_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3002__B _4233_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3768__A2 _3767_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2976__B1 _3669_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2841__B _2841_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput308 _2800_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__3953__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4177_/CLK _4170_/D vssd1 vssd1 vccd1 vccd1 _4170_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3153__A0 _3167_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3391__C _3400_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2900__A0 _3245_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3121_ _3243_/C _4207_/Q _3147_/S vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _3063_/A _3052_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3053_/A sky130_fd_sc_hd__and3_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2003_ input33/X _2001_/X _2002_/Y _1962_/A vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__o211ai_4
XFILLER_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3759__A2 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3954_ _3954_/A vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2967__B1 _3661_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2431__A2 _2428_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3847__B _3853_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2905_ _3861_/A _4035_/Q _2905_/S vssd1 vssd1 vccd1 vccd1 _3247_/C sky130_fd_sc_hd__mux2_2
X_3885_ _3885_/A _3893_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__and3_1
X_2836_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2885_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2767_ _2767_/A _2780_/B _3370_/C vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__and3_2
XANTENNA__3863__A _3871_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2698_ _3291_/C _4121_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3931__A2 _3908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3582__B _3586_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3144__A0 _3262_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2352__D1 _2352_/D1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2498__A2 _3543_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4368_ _4380_/CLK _4368_/D vssd1 vssd1 vccd1 vccd1 _4368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input5_A cpu_adr_i[12] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4346_/CLK _4299_/D vssd1 vssd1 vccd1 vccd1 _4299_/Q sky130_fd_sc_hd__dfxtp_1
X_3319_ _4061_/Q _3314_/X _2165_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _4061_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3998__A2 _3992_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3103__A _3117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4132__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2958__A0 _3798_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4282__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3195__D _3219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__A2 _3902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3492__B _4131_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1933__A1 _1930_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2489__A2 _2485_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3013__A _3021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2110__A1 _2384_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output217_A _3104_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__A _4002_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2852__A _2859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2949__A0 _4288_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3667__B _3796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3159__S _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3386__C _3400_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3670_ _3670_/A vssd1 vssd1 vccd1 vccd1 _4222_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3683__A _3935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2621_ _2427_/A _2428_/A _2517_/X _2434_/A _4386_/Q vssd1 vssd1 vccd1 vccd1 _2621_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2177__A1 _2038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2552_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3913__A2 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput149 _2500_/X vssd1 vssd1 vccd1 vccd1 cpu_dat_o[14] sky130_fd_sc_hd__buf_2
X_2483_ _2382_/X _2383_/X _2483_/C _2503_/D vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__and4bb_1
X_4222_ _4250_/CLK _4222_/D vssd1 vssd1 vccd1 vccd1 _4222_/Q sky130_fd_sc_hd__dfxtp_1
X_4153_ _4389_/CLK _4153_/D vssd1 vssd1 vccd1 vccd1 _4153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2746__B _4142_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3104_ _3104_/A vssd1 vssd1 vccd1 vccd1 _3104_/X sky130_fd_sc_hd__clkbuf_1
X_4084_ _4284_/CLK _4084_/D vssd1 vssd1 vccd1 vccd1 _4084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _3035_/A vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4155__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2762__A _2762_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3858__A _3871_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3937_ _2059_/B _2059_/C _3912_/Y vssd1 vssd1 vccd1 vccd1 _4353_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__3069__S _3076_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3868_ _3868_/A vssd1 vssd1 vccd1 vccd1 _4318_/D sky130_fd_sc_hd__clkbuf_1
X_2819_ _2819_/A vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3593__A _3617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3799_ _3799_/A vssd1 vssd1 vccd1 vccd1 _4290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3904__A2 _3902_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2340__A1 _3530_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A spi_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input80_A gpio_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput18 cpu_adr_i[24] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput29 cpu_adr_i[5] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4028__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3008__A _3010_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output167_A _2642_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2316__D1 _2315_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2847__A _2859_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__CLK _4388_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2331__A1 _2330_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1971__A_N input5/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2634__A2 _2387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2095__B1 _1974_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3678__A _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2582__A _2582_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ _1983_/A _2081_/B _2053_/A _2081_/D vssd1 vssd1 vccd1 vccd1 _1983_/Y sky130_fd_sc_hd__nand4_4
X_3722_ _3722_/A vssd1 vssd1 vccd1 vccd1 _4247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _3653_/A _3661_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__and3_1
X_2604_ _2423_/A _2446_/X _4173_/Q vssd1 vssd1 vccd1 vccd1 _2604_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__1926__A _4357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3584_ _3584_/A _3584_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__and3_1
XFILLER_88_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2535_ _2481_/X _2501_/X _2429_/X _2434_/X _4375_/Q vssd1 vssd1 vccd1 vccd1 _2535_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2570__A1 _2512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2466_ _2507_/A _3677_/A _2507_/C _2466_/D vssd1 vssd1 vccd1 vccd1 _2466_/Y sky130_fd_sc_hd__nand4_1
X_4205_ _4275_/CLK _4205_/D vssd1 vssd1 vccd1 vccd1 _4205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2757__A _2958_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4136_ _4141_/CLK _4136_/D vssd1 vssd1 vccd1 vccd1 _4136_/Q sky130_fd_sc_hd__dfxtp_1
X_2397_ _2390_/Y _3673_/B _2396_/Y vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2476__B _2520_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4302_/CLK _4067_/D vssd1 vssd1 vccd1 vccd1 _4067_/Q sky130_fd_sc_hd__dfxtp_1
X_3018_ _3018_/A vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2625__A2 _2256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2492__A _2590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3588__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2923__C _3431_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2389__A1 _3536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2010__B1 _2009_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2561__A1 _2561_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4320__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2616__A2 _2406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2077__B1 _4069_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3010__B _4237_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3945__B _3965_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3664__C _3664_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output284_A _2842_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3961__A _3961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2320_ _2319_/X _2289_/X _4150_/Q vssd1 vssd1 vccd1 vccd1 _2320_/Y sky130_fd_sc_hd__a21boi_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2644_/A sky130_fd_sc_hd__buf_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__B1 _3489_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2296__B _2393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2182_ _2182_/A _2182_/B vssd1 vssd1 vccd1 vccd1 _2184_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2068__B1 _4072_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3839__C _3839_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3201__A _3201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2462__D _2503_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1966_ _1965_/X _1942_/B _1918_/Y _4285_/Q _4146_/Q vssd1 vssd1 vccd1 vccd1 _1967_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3705_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3855__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2791__A1 _4086_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4343__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3636_ _3636_/A vssd1 vssd1 vccd1 vccd1 _4208_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3574__C _3657_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4389__D _4389_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3567_ _4180_/Q _3523_/X _2407_/X _3566_/X vssd1 vssd1 vccd1 vccd1 _4180_/D sky130_fd_sc_hd__o211a_1
X_2518_ _2363_/X _2449_/X _2517_/X _2450_/X _4374_/Q vssd1 vssd1 vccd1 vccd1 _2518_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3871__A _3871_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3498_ _4134_/Q _3488_/X _3489_/X _3490_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _4134_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2487__A _2507_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2449_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__buf_4
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2310__A4 _2421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4119_ _4251_/CLK _4119_/D vssd1 vssd1 vccd1 vccd1 _4119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3111__A _3111_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3559__B1 _2613_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4299__D _4299_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2534__A1 _4268_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2534__B2 input82/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A cpu_dat_i[17] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2828__C _3394_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4216__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3021__A _3021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3659__C _3659_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2470__B1 _2404_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2860__A _2860_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4366__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3675__B _3796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2222__B1 _2429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3394__C _3394_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__B1 _2417_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3421_ _3421_/A vssd1 vssd1 vccd1 vccd1 _4103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2525__A1 _2512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3352_ _3942_/A _3942_/C _3349_/X _3350_/X _3351_/X vssd1 vssd1 vccd1 vccd1 _4076_/D
+ sky130_fd_sc_hd__o2111a_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2429_/A vssd1 vssd1 vccd1 vccd1 _2303_/X sky130_fd_sc_hd__buf_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3283_ _3320_/A _3283_/B _3323_/C _3317_/C vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__or4_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2234_ _2393_/A vssd1 vssd1 vccd1 vccd1 _2335_/A sky130_fd_sc_hd__clkbuf_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2028_/A _2001_/X _2164_/Y _2184_/C vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ _1965_/X _1942_/B _1918_/Y _4286_/Q _4250_/Q vssd1 vssd1 vccd1 vccd1 _2207_/D
+ sky130_fd_sc_hd__a311oi_2
XANTENNA__3789__B1 _3748_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__C _3657_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2461__B1 _2377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3288__D _3317_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3866__A _3866_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2998_ _2998_/A vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2213__B1 _4217_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1949_ _4057_/Q vssd1 vssd1 vccd1 vccd1 _1949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2764__A1 _4012_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3619_ _3619_/A vssd1 vssd1 vccd1 vccd1 _4200_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3713__B1 _3696_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2516__A1 _2516_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3106__A _3117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4239__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4389__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2680__A _3190_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2504__B1_N _4162_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3942__C _3942_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output247_A _2658_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3016__A _3016_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2691__B1 _3459_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3389__C _3389_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3970_ _3968_/X _3969_/X _2417_/X _2432_/Y vssd1 vssd1 vccd1 vccd1 _4366_/D sky130_fd_sc_hd__o22a_1
XANTENNA__2443__B1 _2404_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2921_ _3867_/C _4038_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _3257_/B sky130_fd_sc_hd__mux2_4
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3686__A _3699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2590__A _2590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2852_ _2859_/A _2872_/B _3402_/C vssd1 vssd1 vccd1 vccd1 _2853_/A sky130_fd_sc_hd__and3_1
XANTENNA__3538__A3 _3528_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2783_ _3447_/B vssd1 vssd1 vccd1 vccd1 _2812_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__1918__B _1923_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3404_ _3444_/A vssd1 vssd1 vccd1 vccd1 _3424_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1934__A _1934_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4384_ _4388_/CLK _4384_/D vssd1 vssd1 vccd1 vccd1 _4384_/Q sky130_fd_sc_hd__dfxtp_1
X_3335_ _3335_/A vssd1 vssd1 vccd1 vccd1 _3724_/D sky130_fd_sc_hd__buf_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3266_ _3266_/A vssd1 vssd1 vccd1 vccd1 _4041_/D sky130_fd_sc_hd__clkbuf_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2197_/X _2200_/X _3052_/B vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2765__A _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _3197_/A vssd1 vssd1 vccd1 vccd1 _3293_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2148_ _4349_/Q _2659_/A _2078_/Y vssd1 vssd1 vccd1 vccd1 _2148_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2682__A0 _3891_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ _4349_/Q _2012_/B _2078_/Y _2137_/A _1985_/X vssd1 vssd1 vccd1 vccd1 _2083_/B
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__3299__C _3323_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3777__A3 _3765_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3596__A _3596_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3529__A3 _3528_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_18_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3934__B1 _2081_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3698__C1 _3683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4061__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2370__C1 _2409_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__A0 _4327_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2976__A1 _2972_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2841__C _3398_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output197_A _3033_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3953__B _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput309 _2807_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3153__A1 _4181_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2900__A1 _4104_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3120_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3147_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _3190_/B _4188_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3586_/C sky130_fd_sc_hd__mux2_1
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2664__A0 _3885_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2002_ _1930_/X _1932_/X _4333_/Q vssd1 vssd1 vccd1 vccd1 _2002_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2967__A1 _2197_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2416__B1 _2415_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3953_ _3953_/A _3953_/B _3953_/C vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__and3_1
XANTENNA__1929__A _4357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3847__C _3847_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2904_ _4315_/Q input51/X _2904_/S vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__mux2_8
XFILLER_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3884_ _3884_/A vssd1 vssd1 vccd1 vccd1 _3914_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2835_ _2835_/A vssd1 vssd1 vccd1 vccd1 _2835_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2766_ _3186_/B _4082_/Q _2937_/S vssd1 vssd1 vccd1 vccd1 _3370_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4084__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3863__B _3877_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2697_ _3898_/A _4051_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _3291_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3582__C _3582_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3144__A1 _4214_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4367_ _4371_/CLK _4367_/D vssd1 vssd1 vccd1 vccd1 _4367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2352__C1 _2286_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3318_ _3318_/A vssd1 vssd1 vccd1 vccd1 _4060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4302_/CLK _4298_/D vssd1 vssd1 vccd1 vccd1 _4298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3249_ _3343_/B vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2655__A0 _3882_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3103__B _3106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3080__A0 _3215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2958__A1 _4010_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3492__C _3502_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1933__A2 _1932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4100__D _4100_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2646__B1 _2298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3013__B _4238_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2110__A2 _2382_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2852__B _2872_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3667__C _3675_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2949__A1 input68/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2620_ _2620_/A1 _2628_/A _2514_/X _2531_/A _2619_/Y vssd1 vssd1 vccd1 vccd1 _3560_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__3964__A _3964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2551_ _4270_/Q _2322_/X _2298_/A input84/X vssd1 vssd1 vccd1 vccd1 _2551_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__2177__A2 _3902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2482_ _2481_/X _2376_/X _2377_/X _2434_/X _4371_/Q vssd1 vssd1 vccd1 vccd1 _2482_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _4225_/CLK _4221_/D vssd1 vssd1 vccd1 vccd1 _4221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3531__D1 _2419_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__D _4010_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4152_ _4388_/CLK _4152_/D vssd1 vssd1 vccd1 vccd1 _4152_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2885__A0 _4312_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _3117_/A _3106_/B _3622_/C vssd1 vssd1 vccd1 vccd1 _3104_/A sky130_fd_sc_hd__and3_1
X_4083_ _4085_/CLK _4083_/D vssd1 vssd1 vccd1 vccd1 _4083_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1931__B _2023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3034_ _3036_/A _4248_/Q vssd1 vssd1 vccd1 vccd1 _3035_/A sky130_fd_sc_hd__and2_1
XANTENNA__2320__B1_N _4150_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3204__A _3224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3858__B _3877_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3062__A0 _3199_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _4352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3867_ _3871_/A _3877_/B _3867_/C vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__or3_1
XANTENNA__3874__A _3874_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2818_ _2828_/A _2841_/B _3389_/C vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__and3_1
X_3798_ _3798_/A _3805_/B _3798_/C vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__or3_1
X_2749_ _2749_/A vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3085__S _3112_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2573__C1 _4380_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2325__C1 _4361_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2876__A0 _3847_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2340__A2 _2255_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3114__A _3114_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A spi_ack_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 cpu_adr_i[25] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input73_A gpio_ack_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2564__C1 _2524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3008__B _4236_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_2_0_CLK_A clkbuf_2_3_0_CLK/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2316__C1 _2409_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2847__B _2872_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2331__A2 _2424_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3024__A _3032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2095__A1 _1968_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _2078_/D vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3694__A _3694_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3721_ _3767_/A _4247_/Q _3721_/C _3724_/D vssd1 vssd1 vccd1 vccd1 _3722_/A sky130_fd_sc_hd__and4_1
X_3652_ _3680_/A vssd1 vssd1 vccd1 vccd1 _3675_/C sky130_fd_sc_hd__buf_2
XANTENNA__2802__S _2825_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3583_ _3583_/A vssd1 vssd1 vccd1 vccd1 _4186_/D sky130_fd_sc_hd__clkbuf_1
X_2603_ _2581_/X _2582_/X _2602_/Y _2579_/X vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1926__B _2201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2103__A _2590_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2534_ _4268_/Q _2295_/X _3771_/A input82/X vssd1 vssd1 vccd1 vccd1 _2534_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__2555__C1 _2524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2465_ _4262_/Q vssd1 vssd1 vccd1 vccd1 _2465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2570__A2 _2513_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2307__C1 _2125_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1942__A _3953_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2396_ _3137_/A _3677_/A _2507_/C _2396_/D vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__nand4_1
X_4204_ _4280_/CLK _4204_/D vssd1 vssd1 vccd1 vccd1 _4204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2858__A0 _3227_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4135_ _4141_/CLK _4135_/D vssd1 vssd1 vccd1 vccd1 _4135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2476__C _2520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3869__A _3869_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4066_ _4326_/CLK _4066_/D vssd1 vssd1 vccd1 vccd1 _4066_/Q sky130_fd_sc_hd__dfxtp_1
X_3017_ _3021_/A _4240_/Q vssd1 vssd1 vccd1 vccd1 _3018_/A sky130_fd_sc_hd__and2_1
XANTENNA__2773__A _2799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2086__A1 _2129_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2492__B _2557_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2389__A2 _2385_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _4339_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2546__C1 _4376_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2010__A1 _4060_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2561__A2 _3369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2849__A0 _4306_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2227__B1_N _2446_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2683__A _2683_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2077__A1 _1993_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3945__C _3945_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3019__A _3021_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4145__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output277_A _2703_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2537__C1 _2536_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2284_/A vssd1 vssd1 vccd1 vccd1 _2421_/A sky130_fd_sc_hd__buf_4
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__B2 _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3501__A1 _4136_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4295__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2296__C _2336_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2181_ _4064_/Q _1977_/X _2180_/Y vssd1 vssd1 vccd1 vccd1 _2186_/C sky130_fd_sc_hd__o21ai_1
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3689__A _3699_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2068__A1 _2055_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1965_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__buf_4
X_3704_ _3704_/A vssd1 vssd1 vccd1 vccd1 _4237_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2240__A1 _2099_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3855__C _3855_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3635_ _3635_/A _3635_/B _3635_/C vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__or3_1
X_3566_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3566_/X sky130_fd_sc_hd__buf_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3497_ _3497_/A vssd1 vssd1 vccd1 vccd1 _4133_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2768__A _2768_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2517_ _2517_/A vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__buf_4
XANTENNA__3871__B _3877_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2448_ _2448_/A1 _2444_/X _2308_/X _2445_/X _2447_/Y vssd1 vssd1 vccd1 vccd1 _3539_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__2487__B _3677_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2379_ _2375_/X _2376_/X _2377_/X _3769_/A _4365_/Q vssd1 vssd1 vccd1 vccd1 _2379_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _4250_/CLK _4118_/D vssd1 vssd1 vccd1 vccd1 _4118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3599__A _3599_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4049_ _4051_/CLK _4049_/D vssd1 vssd1 vccd1 vccd1 _4049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2462__B_N _2383_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4018__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3559__A1 _3559_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4168__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1990__B1 _1989_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2678__A _2678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2534__A2 _2295_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input36_A cpu_dat_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3302__A _3302_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3021__B _4242_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2470__A1 _2461_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2222__A1 _2452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3675__C _3675_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2222__B2 _2552_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3970__A1 _3968_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__B2 _2432_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3972__A _4002_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3420_ _3420_/A _3429_/B _3424_/C vssd1 vssd1 vccd1 vccd1 _3421_/A sky130_fd_sc_hd__and3_1
XFILLER_98_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2525__A2 _2513_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3351_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3351_/X sky130_fd_sc_hd__buf_4
X_2302_ _3730_/B vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__buf_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3282_ _3295_/C vssd1 vssd1 vccd1 vccd1 _3323_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2233_ _2543_/A _2190_/Y _2231_/Y _2232_/Y vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__a31oi_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2164_ _1952_/X _2160_/X _4341_/Q vssd1 vssd1 vccd1 vccd1 _2164_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3789__A1 _4286_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3212__A _3264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2095_ _1968_/Y _2093_/X _1974_/Y _1990_/Y _3301_/A vssd1 vssd1 vccd1 vccd1 _2098_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3789__B2 _3736_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2461__B2 _2434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2461__A1 _2375_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4310__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2997_ _2999_/A _4231_/Q vssd1 vssd1 vccd1 vccd1 _2998_/A sky130_fd_sc_hd__and2_1
XANTENNA__2213__A1 _2129_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1948_ _4059_/Q _2093_/A _1947_/Y vssd1 vssd1 vccd1 vccd1 _2207_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__3882__A _3895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3618_ _3635_/A _3635_/B _3618_/C vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__or3_1
XANTENNA__3713__A1 _4242_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3713__B2 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2516__A2 _2444_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3549_ _3549_/A vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__buf_2
XFILLER_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3106__B _3106_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3122__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2961__A _3115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2900__S _2911_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4103__D _4103_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1963__B1 _1962_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__A _3792_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2201__A _2201_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2140__B1 _4055_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3032__A _3032_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2691__A1 _2677_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4333__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2443__A1 _2435_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2920_ _4318_/Q input54/X _2940_/S vssd1 vssd1 vccd1 vccd1 _3867_/C sky130_fd_sc_hd__mux2_2
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3686__B _4229_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2590__B _2590_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2851_ _3224_/B _4096_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _3402_/C sky130_fd_sc_hd__mux2_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2782_ _2782_/A vssd1 vssd1 vccd1 vccd1 _3447_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1918__C _1924_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__D _4013_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3403_ _3403_/A vssd1 vssd1 vccd1 vccd1 _4096_/D sky130_fd_sc_hd__clkbuf_1
X_4383_ _4389_/CLK _4383_/D vssd1 vssd1 vccd1 vccd1 _4383_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3207__A _3692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3334_ _4068_/Q _3331_/X _3333_/X _3346_/C vssd1 vssd1 vccd1 vccd1 _4068_/D sky130_fd_sc_hd__a211o_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3265_ _3273_/A _3279_/B _3265_/C _3286_/D vssd1 vssd1 vccd1 vccd1 _3266_/A sky130_fd_sc_hd__and4_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3052_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1950__A _2059_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3196_ _3196_/A vssd1 vssd1 vccd1 vccd1 _4016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2147_ _3346_/A _3346_/B _2060_/Y _2064_/Y _2069_/Y vssd1 vssd1 vccd1 vccd1 _2159_/A
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2682__A1 _4048_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ input19/X _2078_/B _2078_/C _2078_/D vssd1 vssd1 vccd1 vccd1 _2078_/Y sky130_fd_sc_hd__nand4b_4
XANTENNA__2781__A _2781_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__A _3895_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3596__B _3609_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3088__S _3109_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2005__B _3303_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__A1 _4351_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__CLK _4280_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3698__B1 _3696_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3117__A _3117_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2021__A _2078_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__B1 _2408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4356__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input138_A spi_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2122__B1 _2121_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2249__C_N _2384_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2673__A1 input27/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2425__A1 _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2976__A2 _2974_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3953__C _3953_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3027__A _3027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__A _2888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2361__B1 _2360_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3050_ _3050_/A vssd1 vssd1 vccd1 vccd1 _3050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2001_ _2001_/A vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3986__B1_N _2554_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2664__A1 _4045_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3697__A _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2416__A1 _2410_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2805__S _2851_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4008__D _4008_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3952_ _3991_/A vssd1 vssd1 vccd1 vccd1 _3952_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2967__A2 _2200_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2903_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2928_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _4324_/D sky130_fd_sc_hd__clkbuf_1
X_2834_ _2859_/A _2841_/B _3396_/A vssd1 vssd1 vccd1 vccd1 _2835_/A sky130_fd_sc_hd__and3_1
XANTENNA__2106__A _2106_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4229__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2765_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2937_/S sky130_fd_sc_hd__buf_2
XANTENNA__1945__A _2007_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3863__C _3863_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2696_ _4331_/Q input31/X _2953_/S vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__mux2_4
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4379__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4366_ _4390_/CLK _4366_/D vssd1 vssd1 vccd1 vccd1 _4366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2565__B1_N _4168_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2352__B1 _2248_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3317_ _3320_/A _3317_/B _3317_/C _3326_/D vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__or4_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4346_/CLK _4297_/D vssd1 vssd1 vccd1 vccd1 _4297_/Q sky130_fd_sc_hd__dfxtp_1
X_3248_ _3248_/A vssd1 vssd1 vccd1 vccd1 _4035_/D sky130_fd_sc_hd__clkbuf_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2655__A1 _4044_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3179_ _3179_/A vssd1 vssd1 vccd1 vccd1 _4009_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3103__C _3622_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3400__A _3400_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3080__A1 _4196_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2040__C1 _2152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2591__B1 _2590_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3540__C1 _3537_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2686__A _2896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2646__A1 _4282_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2110__A3 _2383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2646__B2 input98/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2852__C _3402_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3310__A _3343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ _3551_/A1 _2283_/X _2286_/X _2549_/Y vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2481_ _3730_/A vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ _4250_/CLK _4220_/D vssd1 vssd1 vccd1 vccd1 _4220_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3531__C1 _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _4389_/CLK _4151_/D vssd1 vssd1 vccd1 vccd1 _4151_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2885__A1 input48/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4082_ _4284_/CLK _4082_/D vssd1 vssd1 vccd1 vccd1 _4082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_17_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3102_ _3231_/B _4202_/Q _3109_/S vssd1 vssd1 vccd1 vccd1 _3622_/C sky130_fd_sc_hd__mux2_1
XANTENNA__1931__C _2022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3033_ _3033_/A vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__B _3204_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3858__C _3858_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3220__A _3220_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3062__A1 _4191_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3935_ _3935_/A _3935_/B _3935_/C vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__or3_1
XANTENNA__4051__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3874__B _3893_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3866_ _3866_/A vssd1 vssd1 vccd1 vccd1 _4317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2817_ _3210_/B _4090_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _3389_/C sky130_fd_sc_hd__mux2_1
X_3797_ _3797_/A vssd1 vssd1 vccd1 vccd1 _4289_/D sky130_fd_sc_hd__clkbuf_1
X_2748_ _2748_/A _4143_/Q vssd1 vssd1 vccd1 vccd1 _2749_/A sky130_fd_sc_hd__and2_1
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3770__C1 _3757_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2573__B1 _2517_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4201__D _4201_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2679_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3890__A _3890_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2325__B1 _2324_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2876__A1 _4030_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1918__A_N _4357_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4349_ _4356_/CLK _4349_/D vssd1 vssd1 vccd1 vccd1 _4349_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3130__A _3130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2261__C1 _4358_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3761__C1 _3755_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2564__B1 _2499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input66_A cpu_dat_i[9] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4111__D _4111_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2316__B1 _2408_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2847__C _3400_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3305__A _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3024__B _4243_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2619__A1 _2423_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output222_A _3118_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4074__CLK _4074_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2095__A2 _2093_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3040__A _3044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _3720_/A vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__buf_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _2078_/C vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3651_ _3651_/A vssd1 vssd1 vccd1 vccd1 _4214_/D sky130_fd_sc_hd__clkbuf_1
X_3582_ _3586_/A _3586_/B _3582_/C vssd1 vssd1 vccd1 vccd1 _3583_/A sky130_fd_sc_hd__or3_1
X_2602_ _2281_/X _2599_/Y _2293_/X _2600_/Y _2601_/Y vssd1 vssd1 vccd1 vccd1 _2602_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__1926__C _1994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2533_ _2533_/A vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__buf_2
XANTENNA__2555__B1 _2554_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4021__D _4021_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _3536_/A _2462_/X _2463_/Y vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2307__B1 _2306_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2395_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2507_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4203_ _4275_/CLK _4203_/D vssd1 vssd1 vccd1 vccd1 _4203_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2858__A1 _4097_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1942__B _1942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4134_ _4141_/CLK _4134_/D vssd1 vssd1 vccd1 vccd1 _4134_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3215__A _3224_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2476__D _2476_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _4074_/CLK _4065_/D vssd1 vssd1 vccd1 vccd1 _4065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3016_ _3016_/A vssd1 vssd1 vccd1 vccd1 _3016_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2773__B _2780_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2086__A2 _2106_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3869__B _3869_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2492__C _2590_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3885__A _3885_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3918_ _3918_/A _3942_/B _3940_/C vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__and3_1
X_3849_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3869_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3743__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2546__B1 _2303_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2010__A2 _2093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2561__A3 _2286_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2849__A1 input41/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3125__A _3135_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2964__A _2964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input120_A spi_dat_i[1] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2077__A2 _2018_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2482__C1 _4371_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4106__D _4106_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__A _3795_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2785__A0 _3813_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3945__D _3945_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2204__A _2204_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3019__B _4241_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2537__B1 _2246_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output172_A _2374_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3035__A _3035_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3501__A2 _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2180_ _2044_/A _2001_/X _2179_/Y _1973_/X _2136_/X vssd1 vssd1 vccd1 vccd1 _2180_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2874__A _2903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3689__B _4231_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2068__A2 _2055_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2473__C1 _4370_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4016__D _4016_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1964_ _4076_/Q vssd1 vssd1 vccd1 vccd1 _2055_/A sky130_fd_sc_hd__inv_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2776__A0 _4294_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3703_ _3717_/A _4237_/Q _3703_/C _3711_/D vssd1 vssd1 vccd1 vccd1 _3704_/A sky130_fd_sc_hd__and4_1
XANTENNA__2240__A2 _2964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _4207_/D sky130_fd_sc_hd__clkbuf_1
X_3565_ _3724_/C vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__clkbuf_4
X_3496_ _3510_/A _4133_/Q _3502_/C vssd1 vssd1 vccd1 vccd1 _3497_/A sky130_fd_sc_hd__and3_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2516_ _2516_/A1 _2444_/X _2514_/X _2445_/X _2515_/Y vssd1 vssd1 vccd1 vccd1 _3546_/B
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__3871__C _3871_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2447_ _2330_/X _2446_/X _4157_/Q vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2487__C _2507_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2378_ _2552_/A vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__buf_4
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _4380_/CLK _4117_/D vssd1 vssd1 vccd1 vccd1 _4117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _4302_/CLK _4048_/D vssd1 vssd1 vccd1 vccd1 _4048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3559__A2 _3365_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2024__A _2024_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3716__C1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1990__A1 _4054_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput290 _2879_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input29_A cpu_adr_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2470__A2 _2468_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4112__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2758__A0 _3802_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2222__A2 _3730_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__A2 _3969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4262__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3350_/X sky130_fd_sc_hd__clkbuf_4
X_2301_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__buf_4
XANTENNA__2930__A0 _4320_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3281_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3320_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ _2422_/A _2446_/A _4179_/Q vssd1 vssd1 vccd1 vccd1 _2232_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _4063_/Q _2093_/X _2162_/Y vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2808__S _2844_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _1976_/Y _2184_/C _1986_/Y vssd1 vssd1 vccd1 vccd1 _3301_/A sky130_fd_sc_hd__o21ai_2
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2109__A _4180_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3789__A2 _2200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2461__A2 _2376_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2996_ _2996_/A vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2213__A2 _2112_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1947_ _1939_/Y _2168_/A _1946_/Y _1977_/A vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__1972__A1 _1951_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _3635_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3882__B _3935_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3713__A2 _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3548_ _4164_/Q _3447_/A _3524_/X _2530_/X _3547_/X vssd1 vssd1 vccd1 vccd1 _4164_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2516__A3 _2514_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2921__A0 _3867_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3299__D_N _1990_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3479_ _4126_/Q _3350_/X _4395_/A _3469_/X _3470_/X vssd1 vssd1 vccd1 vccd1 _4126_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3106__C _3624_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3403__A _3403_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3122__B _3125_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4135__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4285__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1963__A1 _1949_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__B _3796_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3313__A _3881_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2140__A1 _2136_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3032__B _4247_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2691__A2 _2680_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output302_A _2774_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2979__A0 _3286_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2443__A2 _2442_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3686__C _3703_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2850_ _3839_/C _4026_/Q _2886_/S vssd1 vssd1 vccd1 vccd1 _3224_/B sky130_fd_sc_hd__mux2_4
XANTENNA__2590__C _2590_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__C1 _3912_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2781_ _2781_/A vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3983__A _3983_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3156__B1 _3572_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3402_ _3407_/A _3413_/B _3402_/C vssd1 vssd1 vccd1 vccd1 _3403_/A sky130_fd_sc_hd__or3_1
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4382_ _4390_/CLK _4382_/D vssd1 vssd1 vccd1 vccd1 _4382_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4008__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3333_ _2201_/X input18/X _1918_/Y _3805_/B _2155_/X vssd1 vssd1 vccd1 vccd1 _3333_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264_ _3264_/A vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4158__CLK _4172_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2215_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__buf_2
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3223__A _3343_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3195_ _3195_/A _3195_/B _3195_/C _3219_/D vssd1 vssd1 vccd1 vccd1 _3196_/A sky130_fd_sc_hd__or4_1
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2146_ _2146_/A _2146_/B _2210_/A vssd1 vssd1 vccd1 vccd1 _2188_/A sky130_fd_sc_hd__nor3_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2077_ _1993_/X _2018_/X _4069_/Q vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__o21ai_1
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3877__B _3877_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3596__C _3600_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2979_ _3286_/C _4223_/Q _3157_/S vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3893__A _3893_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4204__D _4204_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2005__C _2005_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__A2 _3908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2302__A _3730_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3147__A0 _3265_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3698__A1 _4234_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3698__B2 _3697_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3117__B _3125_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2370__A1 _2262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3133__A _3133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2122__A1 _1942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2972__A _3036_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2425__A2 _2424_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input96_A gpio_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4114__D _4114_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2911__S _2911_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3138__A0 _3257_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__A _3308_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2212__A _2964_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output252_A _2716_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2361__A1 _2361_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4300__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__B _2872_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2649__C1 _2648_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _1993_/X _1996_/X _4053_/Q vssd1 vssd1 vccd1 vccd1 _2145_/C sky130_fd_sc_hd__o21ai_1
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3978__A _3978_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3951_ _3728_/A _2260_/X _3945_/D _3800_/A _2380_/A vssd1 vssd1 vccd1 vccd1 _3991_/A
+ sky130_fd_sc_hd__o2111a_2
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2902_ _2902_/A vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2416__A2 _2411_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3882_ _3895_/A _3935_/B _3882_/C vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__or3_1
X_2833_ _3217_/C _4093_/Q _2858_/S vssd1 vssd1 vccd1 vccd1 _3396_/A sky130_fd_sc_hd__mux2_2
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4024__D _4024_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2764_ _3805_/C _4012_/Q _2954_/S vssd1 vssd1 vccd1 vccd1 _3186_/B sky130_fd_sc_hd__mux2_2
XANTENNA__2821__S _2845_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2695_ _2677_/X _2680_/X _3462_/C vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__o21a_2
XANTENNA__3218__A _3218_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4365_ _4371_/CLK _4365_/D vssd1 vssd1 vccd1 vccd1 _4365_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2352__A1 _2700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1961__A _1961_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _4059_/Q _3314_/X _1947_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _4059_/D sky130_fd_sc_hd__o211a_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4302_/CLK _4296_/D vssd1 vssd1 vccd1 vccd1 _4296_/Q sky130_fd_sc_hd__dfxtp_1
X_3247_ _3247_/A _3253_/B _3247_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3248_/A sky130_fd_sc_hd__and4_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3178_ _3192_/A _3199_/B _3178_/C _3945_/A vssd1 vssd1 vccd1 vccd1 _3179_/A sky130_fd_sc_hd__and4_1
XANTENNA__2792__A _2799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2129_ _2129_/A _2129_/B vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3888__A _3888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3400__B _3405_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2591__A1 _2589_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2040__B1 _2038_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4323__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2032__A _4066_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3540__B1 _2463_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2646__A2 _2295_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4109__D _4109_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2906__S _2916_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input11_A cpu_adr_i[18] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3798__A _3798_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3310__B _3326_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2207__A _2207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3038__A _3137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2328_/X _2329_/X _3977_/A _2469_/X vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__o211a_1
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _4172_/CLK _4150_/D vssd1 vssd1 vccd1 vccd1 _4150_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3531__B1 _2356_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3101_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3117_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4081_ _4225_/CLK _4081_/D vssd1 vssd1 vccd1 vccd1 _4081_/Q sky130_fd_sc_hd__dfxtp_1
X_3032_ _3032_/A _4247_/Q vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__and2_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__C _3224_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2816__S _2826_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4019__D _4019_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2117__A _4284_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3934_ _4351_/Q _3908_/A _2081_/Y _3349_/X _3938_/A vssd1 vssd1 vccd1 vccd1 _4351_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3865_ _3865_/A _3869_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__and3_1
X_2816_ _3823_/C _4020_/Q _2826_/S vssd1 vssd1 vccd1 vccd1 _3210_/B sky130_fd_sc_hd__mux2_4
XANTENNA__3874__C _3879_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1956__A _2078_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4346__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3796_ _3796_/A _3796_/B _3903_/A vssd1 vssd1 vccd1 vccd1 _3797_/A sky130_fd_sc_hd__and3_1
X_2747_ _2747_/A vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2678_ _2678_/A vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__buf_4
XANTENNA__2573__B2 _2450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3770__B1 _2558_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2573__A1 _2363_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2787__A _2799_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2325__B2 _2304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2325__A1 _2301_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _4356_/CLK _4348_/D vssd1 vssd1 vccd1 vccd1 _4348_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input3_A cpu_adr_i[10] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4279_ _4286_/CLK _4279_/D vssd1 vssd1 vccd1 vccd1 _4279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A _3411_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2027__A _2027_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2261__B1 _3728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2013__B1 _4342_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3761__B1 _3754_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2564__A1 _2559_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input59_A cpu_dat_i[31] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2316__A1 _2262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2619__A2 _2387_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4219__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output215_A _3097_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3321__A _3321_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3040__B _3052_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4369__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1980_ _2078_/B vssd1 vssd1 vccd1 vccd1 _2081_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3650_ _3659_/A _3659_/B _3650_/C vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__or3_1
X_2601_ _2407_/A _2302_/X _2324_/X _2552_/X _4383_/Q vssd1 vssd1 vccd1 vccd1 _2601_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3581_ _3581_/A vssd1 vssd1 vccd1 vccd1 _4185_/D sky130_fd_sc_hd__clkbuf_1
X_2532_ _3466_/C _4164_/Q _2530_/X _3544_/A vssd1 vssd1 vccd1 vccd1 _2532_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__3991__A _3991_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2555__A1 _2512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4302__D _4302_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2463_ _2287_/X _3468_/A _4158_/Q vssd1 vssd1 vccd1 vccd1 _2463_/Y sky130_fd_sc_hd__a21boi_1
X_4202_ _4280_/CLK _4202_/D vssd1 vssd1 vccd1 vccd1 _4202_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2307__A1 _2224_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2394_ _2638_/B vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2400__A _2474_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1942__C _2023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4133_ _4141_/CLK _4133_/D vssd1 vssd1 vccd1 vccd1 _4133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3215__B _3215_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4064_ _4326_/CLK _4064_/D vssd1 vssd1 vccd1 vccd1 _4064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3015_ _3021_/A _4239_/Q vssd1 vssd1 vccd1 vccd1 _3016_/A sky130_fd_sc_hd__and2_1
XFILLER_97_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2773__C _3372_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3231__A _3250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3869__C _3879_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2492__D _2492_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2048__A_N _2182_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3885__B _3893_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2243__B1 _2239_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3917_ _1939_/Y _3902_/A _1946_/Y vssd1 vssd1 vccd1 vccd1 _3918_/A sky130_fd_sc_hd__o21ai_1
X_3848_ _3848_/A vssd1 vssd1 vccd1 vccd1 _4310_/D sky130_fd_sc_hd__clkbuf_1
X_3779_ _3769_/X _3764_/X _3765_/X _2609_/Y _3774_/X vssd1 vssd1 vccd1 vccd1 _4277_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4212__D _4212_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3743__B1 _2338_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2546__B2 _2304_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2546__A1 _2427_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3406__A _3406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_20_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4225_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3125__B _3125_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input113_A spi_dat_i[13] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__B1 _2377_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2785__A1 _4015_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4122__D _4122_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2537__A1 _2512_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output165_A _2633_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__C1 _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2220__A _2517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_11_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4251_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4041__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3689__C _3703_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4191__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2473__B1 _2311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2890__A _2919_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ _1949_/Y _2184_/C _1962_/Y vssd1 vssd1 vccd1 vccd1 _3308_/C sky130_fd_sc_hd__o21ai_1
X_3702_ _3720_/A vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2776__A1 input60/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3633_ _3633_/A _3633_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__and3_1
XANTENNA__4032__D _4032_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3564_ _3564_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _4179_/D sky130_fd_sc_hd__nor2_1
X_3495_ _3516_/A vssd1 vssd1 vccd1 vccd1 _3510_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2515_ _2330_/X _2446_/X _4163_/Q vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__a21boi_1
X_2446_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2130__A _2130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3226__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2487__D _2487_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4116_ _4250_/CLK _4116_/D vssd1 vssd1 vccd1 vccd1 _4116_/Q sky130_fd_sc_hd__dfxtp_1
X_2377_ _3728_/A vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4047_ _4051_/CLK _4047_/D vssd1 vssd1 vccd1 vccd1 _4047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2464__B1 _2463_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4207__D _4207_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3896__A _3896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3559__A3 _3544_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3716__B1 _3044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2024__B _2072_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1990__A2 _2093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4064__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput280 _2762_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__3136__A _3136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput291 _2768_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_88_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4117__D _4117_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2914__S _2935_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_0_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4356_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2215__A _3054_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2758__A1 _4011_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1966__C1 _4146_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output282_A _2829_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3046__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2300_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2427_/A sky130_fd_sc_hd__buf_4
XANTENNA__2930__A1 input56/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3280_ _3280_/A vssd1 vssd1 vccd1 vccd1 _4047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2678_/A _3269_/C vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__nand2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2143__C1 _3332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2694__A0 _3288_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ _2024_/A _2001_/X _2161_/Y _1973_/X _1965_/X vssd1 vssd1 vccd1 vccd1 _2162_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2093_ _2093_/A vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__buf_2
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4027__D _4027_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2995_ _2999_/A _4230_/Q vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__and2_1
XANTENNA__2125__A _2579_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4087__CLK _4225_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1946_ _2120_/A _2141_/A _4339_/Q vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__1964__A _4076_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3616_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1972__A2 _1994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3882__C _3882_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3547_ _3547_/A vssd1 vssd1 vccd1 vccd1 _3547_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2516__A4 _2445_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2921__A1 _4038_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3478_ _3478_/A vssd1 vssd1 vccd1 vccd1 _4125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2429_ _2429_/A vssd1 vssd1 vccd1 vccd1 _2429_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2685__B1 _3457_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3122__C _3633_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3937__B1 _3912_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2070__D1 _2069_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1963__A2 _2184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__C _3903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A cpu_dat_i[15] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2909__S _2940_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2676__B1 _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2140__A2 _3942_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2979__A1 _4223_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3686__D _3689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2590__D _2590_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__B1 _3927_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2780_ _2799_/A _2780_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _2781_/A sky130_fd_sc_hd__and3_2
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2600__B1 _2298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3156__A1 _2988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4381_ _4389_/CLK _4381_/D vssd1 vssd1 vccd1 vccd1 _4381_/Q sky130_fd_sc_hd__dfxtp_1
X_3401_ _3401_/A vssd1 vssd1 vccd1 vccd1 _4095_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2272__C_N input73/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2364__C1 _4364_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4310__D _4310_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3332_ _3332_/A vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__clkbuf_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3263_ _3263_/A vssd1 vssd1 vccd1 vccd1 _4040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3504__A _3935_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2214_ _2139_/Y _3115_/A _2213_/Y vssd1 vssd1 vccd1 vccd1 _3054_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2667__A0 _3273_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3194_ _3343_/B vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2145_ _3294_/C _3294_/B _2145_/C _2145_/D vssd1 vssd1 vccd1 vccd1 _2210_/A sky130_fd_sc_hd__nand4_1
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2076_ _2076_/A _2076_/B _2158_/C vssd1 vssd1 vccd1 vccd1 _2084_/A sky130_fd_sc_hd__nand3_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3092__A0 _3221_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__C _3877_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1959__A _2023_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2978_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3157_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__3893__B _3893_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1929_ _4357_/Q vssd1 vssd1 vccd1 vccd1 _1951_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2005__D _2098_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3147__A1 _4215_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3698__A2 _3695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4220__D _4220_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3117__C _3631_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2370__A2 _2375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__B1 _3449_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4102__CLK _4180_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3414__A _3414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2122__A2 _1971_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4252__CLK _4284_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input89_A gpio_dat_i[23] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3138__A1 _4212_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__B _3774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4130__D _4130_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2897__A0 _4314_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output245_A _4394_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2361__A2 _2090_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2866__C _3407_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3324__A _3324_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2649__B1 _2469_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3950_ _3950_/A vssd1 vssd1 vccd1 vccd1 _4358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2901_ _2917_/A _2901_/B _3422_/C vssd1 vssd1 vccd1 vccd1 _2902_/A sky130_fd_sc_hd__and3_1
XANTENNA__2821__A0 _3826_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__buf_2
XANTENNA__4305__D _4305_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2081__A_N _2150_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2832_ _3831_/A _4023_/Q _2845_/S vssd1 vssd1 vccd1 vccd1 _3217_/C sky130_fd_sc_hd__mux2_2
X_2763_ _4292_/Q input46/X _2953_/S vssd1 vssd1 vccd1 vccd1 _3805_/C sky130_fd_sc_hd__mux2_1
X_2694_ _3288_/B _4120_/Q _3161_/A vssd1 vssd1 vccd1 vccd1 _3462_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4125__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4040__D _4040_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _4388_/CLK _4364_/D vssd1 vssd1 vccd1 vccd1 _4364_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2352__A2 _2678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3315_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3315_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1961__B _1998_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _4346_/CLK _4295_/D vssd1 vssd1 vccd1 vccd1 _4295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3246_ _3246_/A vssd1 vssd1 vccd1 vccd1 _4034_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3234__A _3247_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4275__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3199_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2128_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2128_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2792__B _2812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _2059_/A _2059_/B _2059_/C vssd1 vssd1 vccd1 vccd1 _2059_/Y sky130_fd_sc_hd__nand3_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3400__C _3400_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4215__D _4215_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2025__D1 _1985_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2313__A _4253_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3409__A _3433_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2040__A1 _4347_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2591__A2 _3617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3540__A1 _2462_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2500__C1 _2469_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3798__B _3805_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3056__A0 _3192_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2803__A0 _3819_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2207__B _2207_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3310__C _3323_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4125__D _4125_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2922__S _2942_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output195_A _3029_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4148__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2223__A _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3531__A1 _2353_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4298__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3100_ _3100_/A vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3054__A _3054_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4080_ _4250_/CLK _4080_/D vssd1 vssd1 vccd1 vccd1 _4080_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3989__A _3989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3031_ _3031_/A vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__D _3219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3933_ input20/X _3908_/X _3932_/X _3912_/Y vssd1 vssd1 vccd1 vccd1 _4350_/D sky130_fd_sc_hd__a211o_1
XANTENNA__4035__D _4035_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3864_ _3864_/A vssd1 vssd1 vccd1 vccd1 _4316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2832__S _2845_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2815_ _4300_/Q input66/X _2825_/S vssd1 vssd1 vccd1 vccd1 _3823_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3229__A _3297_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3795_ _3795_/A vssd1 vssd1 vccd1 vccd1 _4288_/D sky130_fd_sc_hd__clkbuf_1
X_2746_ _2748_/A _4142_/Q vssd1 vssd1 vccd1 vccd1 _2747_/A sky130_fd_sc_hd__and2_1
XANTENNA__2133__A _2133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2677_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3770__A1 _3769_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2573__A2 _2449_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2787__B _2812_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2325__A2 _2302_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _4347_/CLK _4347_/D vssd1 vssd1 vccd1 vccd1 _4347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4278_ _4282_/CLK _4278_/D vssd1 vssd1 vccd1 vccd1 _4278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3229_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3250_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3899__A _3899_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2494__D1 _2493_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2308__A _2514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2261__A1 _2256_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2261__B2 _2260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3139__A _3151_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2043__A _2043_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2013__A1 _1930_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3761__A1 _4266_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3761__B2 _2507_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2978__A _3206_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2564__A2 _2563_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2316__A2 _2375_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3602__A _3611_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output208_A _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2218__A _2346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3040__C _3580_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2652__S _2949_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3049__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2600_ _4276_/Q _2322_/X _2298_/A input91/X vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__a22oi_4
X_3580_ _3580_/A _3584_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3581_/A sky130_fd_sc_hd__and3_1
X_2531_ _2531_/A vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2888__A _2888_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2555__A2 _2513_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2462_ _2382_/X _2383_/X _2462_/C _2503_/D vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__2307__A2 _2245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4201_ _4201_/CLK _4201_/D vssd1 vssd1 vccd1 vccd1 _4201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2393_ _2393_/A vssd1 vssd1 vccd1 vccd1 _2638_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1942__D _2022_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _4177_/CLK _4132_/D vssd1 vssd1 vccd1 vccd1 _4132_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3215__C _3224_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2827__S _2851_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4063_ _4326_/CLK _4063_/D vssd1 vssd1 vccd1 vccd1 _4063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _3014_/A vssd1 vssd1 vccd1 vccd1 _3014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3231__B _3231_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2128__A _2752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4313__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2243__A1 _2418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1967__A _2207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3885__C _3914_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3916_ _3938_/A _3916_/B _3916_/C _3938_/D vssd1 vssd1 vccd1 vccd1 _4338_/D sky130_fd_sc_hd__nand4_1
XANTENNA__2243__B2 _2292_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3847_ _3847_/A _3853_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__or3_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _4276_/Q _3767_/X _3771_/X input91/X _3772_/X vssd1 vssd1 vccd1 vccd1 _4276_/D
+ sky130_fd_sc_hd__a221o_1
X_2729_ _2737_/A _4134_/Q vssd1 vssd1 vccd1 vccd1 _2730_/A sky130_fd_sc_hd__and2_1
XANTENNA__3743__A1 _3727_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2546__A2 _2428_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3125__C _3635_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3422__A _3431_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__B2 _2434_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2482__A1 _2481_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__A _2038_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input106_A gpio_err_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2537__A2 _2513_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input71_A cpu_stb_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2501__A _3730_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3498__B1 _3489_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output158_A _2580_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2170__B1 _2169_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4336__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3332__A _3332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3689__D _3689_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__D1 _2457_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2473__B2 _2450_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2473__A1 _2363_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ _1962_/A _1962_/B _1962_/C vssd1 vssd1 vccd1 vccd1 _1962_/Y sky130_fd_sc_hd__nand3_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3701_ _4236_/Q _3695_/X _3696_/X _3697_/X _3683_/X vssd1 vssd1 vccd1 vccd1 _4236_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3632_ _3632_/A vssd1 vssd1 vccd1 vccd1 _4206_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4313__D _4313_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3507__A _3510_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3563_ _4178_/Q _3447_/A _3524_/X _2644_/X _3549_/A vssd1 vssd1 vccd1 vccd1 _4178_/D
+ sky130_fd_sc_hd__a221o_1
X_3494_ _4132_/Q _3488_/X _3489_/X _3490_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _4132_/D
+ sky130_fd_sc_hd__a221o_1
X_2514_ _2514_/A vssd1 vssd1 vccd1 vccd1 _2514_/X sky130_fd_sc_hd__buf_4
XANTENNA__2411__A _3641_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2445_ _2531_/A vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__buf_4
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2376_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__buf_2
X_4115_ _4251_/CLK _4115_/D vssd1 vssd1 vccd1 vccd1 _4115_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2161__B1 _4343_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3242__A _3242_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4046_ _4085_/CLK _4046_/D vssd1 vssd1 vccd1 vccd1 _4046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2464__A1 _3536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3984__B1_N _2536_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2503__B_N _2383_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4223__D _4223_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1975__B1 _1974_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3716__B2 _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3716__A1 _4244_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4209__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2024__C _2081_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3417__A _3441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput270 _2751_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[30] sky130_fd_sc_hd__buf_2
Xoutput292 _2884_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput281 _2824_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_88_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4359__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3152__A _3152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2991__A _2999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4133__D _4133_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2930__S _2940_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1966__B1 _4285_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output275_A _2695_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3327__A _3327_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2231__A _2678_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _3942_/C _1996_/X _3879_/A _2138_/X vssd1 vssd1 vccd1 vccd1 _3269_/C sky130_fd_sc_hd__o31a_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3340__C1 _3805_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2143__B1 _2142_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2694__A1 _4120_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _1952_/X _2160_/X _4343_/Q vssd1 vssd1 vccd1 vccd1 _2161_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2092_ _2207_/A _2207_/B vssd1 vssd1 vccd1 vccd1 _2098_/A sky130_fd_sc_hd__and2_1
XFILLER_93_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3997__A _3997_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4308__D _4308_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2994_ _2994_/A vssd1 vssd1 vccd1 vccd1 _2994_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2406__A _2406_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _2007_/A vssd1 vssd1 vccd1 vccd1 _2141_/A sky130_fd_sc_hd__buf_2
XANTENNA__2840__S _2851_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4043__D _4043_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3615_ _3615_/A vssd1 vssd1 vccd1 vccd1 _4199_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3237__A _3237_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3546_ _3546_/A _3546_/B vssd1 vssd1 vccd1 vccd1 _4163_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2141__A _2141_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3477_ _3492_/A _4125_/Q _4002_/B vssd1 vssd1 vccd1 vccd1 _3478_/A sky130_fd_sc_hd__and3_1
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1980__A _2078_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2428_ _2428_/A vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__buf_2
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2685__A1 _2677_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2359_ _2328_/X _2329_/X _2246_/X _2358_/Y vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__o211a_1
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2437__A1 _2287_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4218__D _4218_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_15_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4029_ _4199_/CLK _4029_/D vssd1 vssd1 vccd1 vccd1 _4029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3700__A _3700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4031__CLK _4199_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3937__A1 _2059_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1948__B1 _1947_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2070__C1 _2064_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4181__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2051__A _3326_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2986__A _2988_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2676__A1 _2128_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3322__C1 _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input34_A cpu_cyc_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__D _4128_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2925__S _2935_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3610__A _3610_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2226__A _2226_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3928__A1 input16/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2600__A1 _4276_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2600__B2 input91/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3156__A2 _2200_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3057__A _3063_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4380_ _4380_/CLK _4380_/D vssd1 vssd1 vccd1 vccd1 _4380_/Q sky130_fd_sc_hd__dfxtp_1
X_3400_ _3400_/A _3405_/B _3400_/C vssd1 vssd1 vccd1 vccd1 _3401_/A sky130_fd_sc_hd__and3_1
XANTENNA__3561__C1 _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2364__B1 _2311_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3331_ _3940_/C vssd1 vssd1 vccd1 vccd1 _3331_/X sky130_fd_sc_hd__buf_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2896__A _2896_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__B1 _2115_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3262_ _3276_/A _3262_/B _3276_/C _3271_/D vssd1 vssd1 vccd1 vccd1 _3263_/A sky130_fd_sc_hd__or4_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2129_/B _2112_/B _4217_/Q vssd1 vssd1 vccd1 vccd1 _2213_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2667__A1 _4115_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3193_ _3193_/A vssd1 vssd1 vccd1 vccd1 _4015_/D sky130_fd_sc_hd__clkbuf_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2144_ _2140_/Y _2143_/X _1990_/Y _3303_/B vssd1 vssd1 vccd1 vccd1 _2146_/A sky130_fd_sc_hd__o211ai_1
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4038__D _4038_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3520__A _3547_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2075_ _4350_/Q _2012_/B _2074_/Y _1938_/A vssd1 vssd1 vccd1 vccd1 _2158_/C sky130_fd_sc_hd__o211ai_4
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3092__A1 _4199_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4054__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2136__A _2136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2977_ _3115_/A vssd1 vssd1 vccd1 vccd1 _3206_/A sky130_fd_sc_hd__clkbuf_2
X_1928_ input7/X _1970_/A vssd1 vssd1 vccd1 vccd1 _3916_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3893__C _3914_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2355__B1 _2644_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3529_ _3529_/A1 _3523_/X _3528_/X _2320_/Y _3562_/A vssd1 vssd1 vccd1 vccd1 _4150_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__A1 _2128_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2122__A3 _1971_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3430__A _3430_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2594__B1 _2593_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__C _3308_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3605__A _3605_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2897__A1 input50/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2361__A3 _2308_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2649__A1 _2328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output238_A _3068_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4077__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2655__S _2950_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2900_ _3245_/B _4104_/Q _2911_/S vssd1 vssd1 vccd1 vccd1 _3422_/C sky130_fd_sc_hd__mux2_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _3880_/A vssd1 vssd1 vccd1 vccd1 _4323_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2821__A1 _4021_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2831_ _4303_/Q input38/X _2844_/S vssd1 vssd1 vccd1 vccd1 _3831_/A sky130_fd_sc_hd__mux2_8
X_2762_ _2762_/A vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2034__C1 _1938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__B1 _2298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4321__D _4321_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2693_ _3895_/C _4050_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _3288_/B sky130_fd_sc_hd__mux2_4
XFILLER_99_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ _4391_/CLK _4363_/D vssd1 vssd1 vccd1 vccd1 _4363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3314_ _3314_/A vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__buf_2
XANTENNA__1961__C _1971_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _4302_/CLK _4294_/D vssd1 vssd1 vccd1 vccd1 _4294_/Q sky130_fd_sc_hd__dfxtp_1
X_3245_ _3250_/A _3245_/B _3250_/C _3245_/D vssd1 vssd1 vccd1 vccd1 _3246_/A sky130_fd_sc_hd__or4_1
XANTENNA__3234__B _3253_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3176_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__buf_4
X_2127_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2752_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2792__C _3378_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3250__A _3250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ _1952_/A _2160_/A _4353_/Q vssd1 vssd1 vccd1 vccd1 _2059_/C sky130_fd_sc_hd__o21ai_1
XFILLER_54_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2025__C1 _2015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2576__B1 _2575_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4231__D _4231_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2040__A2 _2012_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3540__A2 _3536_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3425__A _3425_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input136_A spi_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2500__B1 _2499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3798__C _3798_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3056__A1 _4189_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2803__A1 _4018_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2207__C _2207_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4005__B1 _2224_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2567__B1 _2298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output188_A _3014_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4141__D _4141_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3531__A2 _3523_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3335__A _3335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3030_ _3032_/A _4246_/Q vssd1 vssd1 vccd1 vccd1 _3031_/A sky130_fd_sc_hd__and2_1
XFILLER_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3989__B _3999_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3070__A _3081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4316__D _4316_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _2121_/X _2201_/X _1994_/X _4350_/Q vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ _3871_/A _3877_/B _3863_/C vssd1 vssd1 vccd1 vccd1 _3864_/A sky130_fd_sc_hd__or3_1
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2814_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2841_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2414__A _2414_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2558__B1 _2557_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3794_ _3798_/A _3805_/B _3794_/C vssd1 vssd1 vccd1 vccd1 _3795_/A sky130_fd_sc_hd__or3_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2745_ _2745_/A vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4051__D _4051_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2676_ _2128_/X _2133_/X _3455_/A vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3770__A2 _3764_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4242__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2787__C _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3245__A _3250_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4346_ _4346_/CLK _4346_/D vssd1 vssd1 vccd1 vccd1 _4346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4280_/CLK _4277_/D vssd1 vssd1 vccd1 vccd1 _4277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3228_ _3228_/A vssd1 vssd1 vccd1 vccd1 _4027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _3180_/B _4184_/Q _3206_/A vssd1 vssd1 vccd1 vccd1 _3576_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2494__C1 _2409_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4226__D _4226_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2797__A0 _3817_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2261__A2 _2258_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2324__A _2429_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3139__B _3142_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3746__C1 _3738_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2013__A2 _1932_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3761__A2 _3750_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2994__A _2994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3602__B _3611_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4136__D _4136_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4115__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2234__A _2393_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3049__B _3052_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2888__B _2901_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2530_ _2628_/A _2644_/B _2530_/C vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__and3_1
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2960__B1 _3365_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2461_ _2375_/X _2376_/X _2377_/X _2434_/X _4369_/Q vssd1 vssd1 vccd1 vccd1 _2461_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3065__A _3696_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4200_ _4280_/CLK _4200_/D vssd1 vssd1 vccd1 vccd1 _4200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2392_ _2412_/A vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__buf_2
X_4131_ _4177_/CLK _4131_/D vssd1 vssd1 vccd1 vccd1 _4131_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3215__D _3219_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4062_ _4326_/CLK _4062_/D vssd1 vssd1 vccd1 vccd1 _4062_/Q sky130_fd_sc_hd__dfxtp_1
X_3013_ _3021_/A _4238_/Q vssd1 vssd1 vccd1 vccd1 _3014_/A sky130_fd_sc_hd__and2_1
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2409__A _2409_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3231__C _3250_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4046__D _4046_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2779__A0 _3190_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1967__B _2207_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _4337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2243__A2 _3564_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3846_ _3846_/A vssd1 vssd1 vccd1 vccd1 _4309_/D sky130_fd_sc_hd__clkbuf_1
X_3777_ _3769_/X _3764_/X _3765_/X _2591_/Y _3774_/X vssd1 vssd1 vccd1 vccd1 _4275_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__1983__A _1983_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2728_ _2739_/A vssd1 vssd1 vccd1 vccd1 _2737_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3743__A2 _3729_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2951__A0 _3174_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2659_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2957_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4346_/CLK _4329_/D vssd1 vssd1 vccd1 vccd1 _4329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3703__A _3717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3422__B _3437_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2319__A _2529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4138__CLK _4141_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1931__A_N _4356_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__A2 _2376_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__B _2072_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3967__C1 _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4288__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2989__A _2989_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3719__C1 _3705_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2942__A0 _3267_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A cpu_dat_i[7] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3498__A1 _4134_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3498__B2 _3490_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3613__A _3666_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2170__A1 _4062_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output220_A _3045_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2458__C1 _2454_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2473__A2 _2449_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _3700_/A vssd1 vssd1 vccd1 vccd1 _4235_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _1961_/A _1998_/B _1971_/C _1971_/D vssd1 vssd1 vccd1 vccd1 _1962_/C sky130_fd_sc_hd__nand4_2
X_3631_ _3635_/A _3635_/B _3631_/C vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__or3_1
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _4177_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3507__B _4139_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2513_ _2582_/A vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3493_ _3493_/A vssd1 vssd1 vccd1 vccd1 _4131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2444_ _2529_/A vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__buf_4
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2375_ _2375_/A vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3523__A _3536_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4114_ _4141_/CLK _4114_/D vssd1 vssd1 vccd1 vccd1 _4114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2161__A1 _1952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4045_ _4199_/CLK _4045_/D vssd1 vssd1 vccd1 vccd1 _4045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2464__A2 _2462_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1978__A _2011_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2621__C1 _4386_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1975__A1 _1968_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3829_ _3847_/A _3829_/B _3829_/C vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__or3_1
XANTENNA__3716__A2 _3167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2024__D _2074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput260 _2732_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput271 _2753_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[31] sky130_fd_sc_hd__buf_2
XFILLER_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput293 _2889_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput282 _2829_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3433__A _3433_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2049__A _2152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2991__B _4228_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2612__C1 _2579_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1966__A1 _1965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3608__A _3608_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2512__A _2581_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2915__A0 _3865_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output268_A _2749_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2231__B _3269_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output170_A _2341_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4303__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__A _3343_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3340__B1 _2074_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2143__A1 _2121_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2160_ _2160_/A vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2091_ _3489_/A vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__buf_2
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2993_ _2999_/A _4229_/Q vssd1 vssd1 vccd1 vccd1 _2994_/A sky130_fd_sc_hd__and2_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2603__C1 _2579_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1944_ _1951_/A vssd1 vssd1 vccd1 vccd1 _2120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4324__D _4324_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3159__A0 _3180_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3614_ _3614_/A _3633_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3615_/A sky130_fd_sc_hd__and3_1
XANTENNA__2422__A _2422_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2906__A0 _3247_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3545_ _2503_/C _3536_/X _3544_/X _2504_/Y _3537_/X vssd1 vssd1 vccd1 vccd1 _4162_/D
+ sky130_fd_sc_hd__a311o_1
X_3476_ _4124_/Q _3350_/X _4395_/A _3469_/X _3470_/X vssd1 vssd1 vccd1 vccd1 _4124_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2427_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__buf_2
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3253__A _3273_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2685__A2 _2680_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2358_ _2342_/Y _2357_/A _2357_/Y vssd1 vssd1 vccd1 vccd1 _2358_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ _2387_/A vssd1 vssd1 vccd1 vccd1 _2289_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4028_ _4380_/CLK _4028_/D vssd1 vssd1 vccd1 vccd1 _4028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2437__A2 _3468_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4234__D _4234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3937__A2 _2059_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2070__B1 _2060_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1948__A1 _4059_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3428__A _3428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4326__CLK _4326_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2051__B _3328_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2986__B _4226_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3163__A _3335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3322__B1 _2162_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2676__A2 _2133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A cpu_adr_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2507__A _2507_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3102__S _3109_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4144__D _4144_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2941__S _2941_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__A2 _3908_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2600__A2 _2322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2005__A_N _2146_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3057__B _3070_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3561__B1 _3524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2364__A1 _2363_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2364__B2 _2260_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3330_ _3790_/A vssd1 vssd1 vccd1 vccd1 _3940_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__A1 input73/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3261_ _3261_/A vssd1 vssd1 vccd1 vccd1 _4039_/D sky130_fd_sc_hd__clkbuf_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3998__B1_N _2617_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2212_ _2964_/A vssd1 vssd1 vccd1 vccd1 _3115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3192_ _3192_/A _3199_/B _3192_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__and4_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4319__D _4319_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2143_ _2121_/X _1983_/A _3953_/B _2142_/Y _3332_/A vssd1 vssd1 vccd1 vccd1 _2143_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3801__A _3897_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ input20/X _2081_/B _2081_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2074_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2851__S _2851_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4349__CLK _4356_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4054__D _4054_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2976_ _2972_/X _2974_/X _3669_/C vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3248__A _3248_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1927_ _2011_/A vssd1 vssd1 vccd1 vccd1 _1970_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2152__A _2152_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2355__A1 _4180_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2355__B2 _2644_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3528_ _3544_/A vssd1 vssd1 vccd1 vccd1 _3528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3459_ _3459_/A _3459_/B _3466_/C vssd1 vssd1 vccd1 vccd1 _3460_/A sky130_fd_sc_hd__and3_1
XANTENNA__2107__A1 _2129_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2658__A2 _2133_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4229__D _4229_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3711__A _3717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2515__B1_N _4163_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2291__B1 _2290_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2594__A1 _2594_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2997__A _2999_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2361__A4 _2421_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3605__B _3609_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4139__D _4139_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2649__A2 _2329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2936__S _2936_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3621__A _3621_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output300_A _2929_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2237__A _2237_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2671__S _2942_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2830_ _3489_/A vssd1 vssd1 vccd1 vccd1 _2859_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ _2767_/A _2780_/B _3367_/A vssd1 vssd1 vccd1 vccd1 _2762_/A sky130_fd_sc_hd__and3_2
XANTENNA__3068__A _3068_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2034__B1 _2033_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__A1 _4274_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__B1 _3771_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__B2 input89/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2692_ _4330_/Q input30/X _2949_/S vssd1 vssd1 vccd1 vccd1 _3895_/C sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_14_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2700__A _2700_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4362_ _4390_/CLK _4362_/D vssd1 vssd1 vccd1 vccd1 _4362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3313_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3314_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1961__D _1971_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4346_/CLK _4293_/D vssd1 vssd1 vccd1 vccd1 _4293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3244_ _3244_/A vssd1 vssd1 vccd1 vccd1 _4033_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3234__C _3234_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2846__S _2858_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4049__D _4049_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3175_ _3175_/A vssd1 vssd1 vccd1 vccd1 _4008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2126_ _4146_/Q vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__buf_2
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4171__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3250__B _3250_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2057_ _2078_/C _2078_/D _2057_/C _2078_/B vssd1 vssd1 vccd1 vccd1 _2059_/B sky130_fd_sc_hd__nand4_2
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2959_ _3180_/B _4080_/Q _3161_/A vssd1 vssd1 vccd1 vccd1 _3365_/C sky130_fd_sc_hd__mux2_4
XANTENNA__2025__B1 _2024_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__B1 _3771_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2576__A1 _2574_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3540__A3 _3528_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2756__S _3907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3441__A _3441_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2500__A1 _2494_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input129_A spi_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2057__A _2078_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2207__D _2207_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4005__B2 _2245_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4005__A1 _3991_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input94_A gpio_dat_i[28] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2016__B1 _4062_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2567__A1 _4272_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2567__B2 input87/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3616__A _3804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2520__A _2575_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4044__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output250_A _2712_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4194__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3989__C _3996_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3351__A _3695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3070__B _3070_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _4349_/Q _3908_/A _2078_/Y _3909_/X _3938_/A vssd1 vssd1 vccd1 vccd1 _4349_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _3862_/A vssd1 vssd1 vccd1 vccd1 _4315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2813_ _2813_/A vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2558__A1 _2556_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4332__D _4332_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3793_ _3793_/A vssd1 vssd1 vccd1 vccd1 _4287_/D sky130_fd_sc_hd__clkbuf_1
X_2744_ _2748_/A _4141_/Q vssd1 vssd1 vccd1 vccd1 _2745_/A sky130_fd_sc_hd__and2_1
XANTENNA__3770__A3 _3765_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2675_ _3279_/C _4117_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__mux2_4
XANTENNA__2430__A _2434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3245__B _3245_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4345_ _4347_/CLK _4345_/D vssd1 vssd1 vccd1 vccd1 _4345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _4282_/CLK _4276_/D vssd1 vssd1 vccd1 vccd1 _4276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3261__A _3261_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3227_ _3247_/A _3227_/B _3227_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _3228_/A sky130_fd_sc_hd__and4_1
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3158_ _2988_/A _2200_/A _3574_/A vssd1 vssd1 vccd1 vccd1 _3158_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2494__B1 _2408_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3691__C1 _3683_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2109_ _4180_/Q vssd1 vssd1 vccd1 vccd1 _2109_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3089_ _3099_/A _3089_/B _3611_/C vssd1 vssd1 vccd1 vccd1 _3090_/A sky130_fd_sc_hd__and3_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3994__B1 _2592_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2797__A1 _4017_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2549__A1 _2319_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4242__D _4242_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3746__B1 _3735_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3139__C _3646_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4067__CLK _4302_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3436__A _3461_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_23_CLK _4201_/CLK vssd1 vssd1 vccd1 vccd1 _4302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3171__A _3591_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2485__B1 _2484_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3602__C _3602_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__B1 _2542_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2331__B1_N _4151_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output298_A _2918_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4152__D _4152_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3737__B1 _3264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3049__C _3584_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4262_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2960__A1 _2704_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2250__A _2284_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2888__C _3418_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2460_ _2328_/X _2329_/X _3973_/A _2373_/X vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3346__A _3346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4130_ _4177_/CLK _4130_/D vssd1 vssd1 vccd1 vccd1 _4130_/Q sky130_fd_sc_hd__dfxtp_1
X_2391_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2173__C1 _2153_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3081__A _3081_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _4326_/CLK _4061_/D vssd1 vssd1 vccd1 vccd1 _4061_/Q sky130_fd_sc_hd__dfxtp_1
X_3012_ _3023_/A vssd1 vssd1 vccd1 vccd1 _3021_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4327__D _4327_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3231__D _3245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2228__B1 _3945_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2779__A1 _4084_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3914_ _3914_/A _3942_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__and3_1
XANTENNA__1967__C _3308_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3845_ _3845_/A _3845_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__and3_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4062__D _4062_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3776_ _4274_/Q _3767_/X _3771_/X input89/X _3772_/X vssd1 vssd1 vccd1 vccd1 _4274_/D
+ sky130_fd_sc_hd__a221o_1
X_2727_ _2727_/A vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3743__A3 _3732_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1983__B _2081_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2951__A1 _4078_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3256__A _3295_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2160__A _2160_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2658_ _2128_/X _2133_/X _3449_/C vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__o21a_1
X_2589_ _4275_/Q vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__B1 _4332_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4328_ _4347_/CLK _4328_/D vssd1 vssd1 vccd1 vccd1 _4328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3703__B _4237_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4259_ _4284_/CLK _4259_/D vssd1 vssd1 vccd1 vccd1 _4259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A RST_N vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3422__C _3422_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4237__D _4237_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2467__B1 _2466_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__C _2081_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2335__A _2335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3967__B1 _2399_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3719__B1 _3044_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2942__A1 _4112_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3166__A _3707_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3498__A2 _3488_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input57_A cpu_dat_i[2] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3352__D1 _3351_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2170__A2 _1977_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3105__S _3112_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4147__D _4147_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2458__B1 _2453_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output213_A _3090_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4232__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4380_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2245__A _2329_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ _2078_/D vssd1 vssd1 vccd1 vccd1 _1971_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2630__B1 _2298_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4382__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3630_ _3630_/A vssd1 vssd1 vccd1 vccd1 _4205_/D sky130_fd_sc_hd__clkbuf_1
X_3561_ _4176_/Q _3447_/A _3524_/X _2628_/X _3549_/A vssd1 vssd1 vccd1 vccd1 _4176_/D
+ sky130_fd_sc_hd__a221o_1
X_2512_ _2581_/A vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3507__C _3657_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3492_ _3492_/A _4131_/Q _3502_/C vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__and3_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2443_ _2435_/X _2442_/Y _2404_/X _2373_/X vssd1 vssd1 vccd1 vccd1 _2443_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3804__A _3804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2374_ _2328_/X _2329_/X _3963_/A _2373_/X vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__o211a_2
XANTENNA__2697__A0 _3898_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4113_ _4180_/CLK _4113_/D vssd1 vssd1 vccd1 vccd1 _4113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2161__A2 _2160_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4085_/CLK _4044_/D vssd1 vssd1 vccd1 vccd1 _4044_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4057__D _4057_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2621__B1 _2517_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1994__A _1994_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3828_ _3876_/A vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1975__A2 _3332_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ _4264_/Q _3750_/X _3754_/X _2487_/D _3755_/X vssd1 vssd1 vccd1 vccd1 _4264_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput261 _2734_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput250 _2712_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__4105__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput272 _2676_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput294 _2895_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput283 _2835_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__3714__A _3717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4255__CLK _4286_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2049__B _3925_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2764__S _2954_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input111_A spi_dat_i[11] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2065__A _2065_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2612__B1 _3996_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2073__D1 _1985_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1966__A2 _1942_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2915__A1 _4037_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output163_A _2618_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3624__A _3624_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3343__B _3343_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3340__A1 _4350_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2143__A2 _1983_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2090_ _2090_/A vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2674__S _2936_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2851__A0 _3224_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2992_ _2992_/A vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2603__B1 _2602_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ _2001_/A vssd1 vssd1 vccd1 vccd1 _2168_/A sky130_fd_sc_hd__buf_2
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2703__A _2703_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3159__A1 _4184_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3613_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3633_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4128__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2906__A1 _4105_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4340__D _4340_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3544_ _3544_/A vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__clkbuf_2
X_3475_ _3475_/A vssd1 vssd1 vccd1 vccd1 _4123_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2849__S _2885_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2426_ _2426_/A1 _2420_/X _2421_/X _2425_/Y vssd1 vssd1 vccd1 vccd1 _3535_/B sky130_fd_sc_hd__a31oi_2
XANTENNA__3534__A _3549_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4278__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3253__B _3253_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2357_ _2357_/A _2357_/B _2357_/C vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__nand3_2
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2288_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2387_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3095__A0 _3224_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4027_ _4199_/CLK _4027_/D vssd1 vssd1 vccd1 vccd1 _4027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3709__A _3709_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2070__A1 _3346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__1948__A2 _2093_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4250__D _4250_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2051__C _2051_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3444__A _3444_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3322__A1 _4063_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2833__A0 _3217_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2507__B _2557_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3619__A _3619_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2597__C1 _2579_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3338__B _3488_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4160__D _4160_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output280_A _2762_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3057__C _3589_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3561__A1 _4176_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3561__B2 _2628_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2364__A2 _2258_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2669__S _2949_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3354__A _3354_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__A2 _2272_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3260_ _3273_/A _3279_/B _3260_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3261_/A sky130_fd_sc_hd__and4_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3191_/A vssd1 vssd1 vccd1 vccd1 _4014_/D sky130_fd_sc_hd__clkbuf_1
X_2211_ _2211_/A _2211_/B _2211_/C _2211_/D vssd1 vssd1 vccd1 vccd1 _2964_/A sky130_fd_sc_hd__nand4_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2142_ _2121_/A _3953_/B _4335_/Q vssd1 vssd1 vccd1 vccd1 _2142_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ _4348_/Q _2012_/B _2072_/Y _2137_/A _1985_/X vssd1 vssd1 vccd1 vccd1 _2076_/B
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4335__D _4335_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2975_ _3283_/B _4222_/Q _3150_/S vssd1 vssd1 vccd1 vccd1 _3669_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2588__C1 _2587_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2052__A1 _2136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1926_ _4357_/Q _2201_/A _1994_/A vssd1 vssd1 vccd1 vccd1 _2011_/A sky130_fd_sc_hd__nor3_1
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4070__D _4070_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3527_ _3564_/B _3527_/B vssd1 vssd1 vccd1 vccd1 _4149_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2355__A2 _2353_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3264__A _3264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3458_ _3458_/A vssd1 vssd1 vccd1 vccd1 _4118_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2107__A2 _2129_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3389_ _3407_/A _3389_/B _3389_/C vssd1 vssd1 vccd1 vccd1 _3390_/A sky130_fd_sc_hd__or3_1
X_2409_ _2409_/A vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3711__B _4241_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2608__A _2638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2815__A0 _4300_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4245__D _4245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2291__A1 _3526_/A1 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__A _3439_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2343__A _4256_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2594__A2 _3369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2997__B _4231_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3174__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3605__C _3624_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3902__A _3902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3059__A0 _3195_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4155__D _4155_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3349__A _3724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2760_ _3184_/C _4081_/Q _2955_/S vssd1 vssd1 vccd1 vccd1 _3367_/A sky130_fd_sc_hd__mux2_2
XANTENNA__2034__A1 input16/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2691_ _2677_/X _2680_/X _3459_/A vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__o21a_2
XANTENNA__3782__A1 _4280_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__A2 _2295_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__B2 input95/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4390_/CLK _4361_/D vssd1 vssd1 vccd1 vccd1 _4361_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3084__A _3120_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3312_ _3332_/A vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__buf_2
X_4292_ _4302_/CLK _4292_/D vssd1 vssd1 vccd1 vccd1 _4292_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3243_ _3247_/A _3253_/B _3243_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3244_/A sky130_fd_sc_hd__and4_1
XANTENNA__3234__D _3234_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3812__A _3884_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3174_ _3195_/A _3174_/B _3195_/C _3190_/D vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__or4_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2428__A _2428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2125_ _2579_/A vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4316__CLK _4391_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3250__C _3250_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2056_ _3938_/B _3938_/C _2134_/A vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__a21oi_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2862__S _2885_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4065__D _4065_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3259__A _3692_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2958_ _3798_/C _4010_/Q _2958_/S vssd1 vssd1 vccd1 vccd1 _3180_/B sky130_fd_sc_hd__mux2_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2025__A1 _4343_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 _4272_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__B2 input87/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2576__A2 _2366_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2889_ _2889_/A vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__A _3722_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2500__A2 _2498_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2057__B _2078_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2772__S _2955_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4005__A2 _3992_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3169__A input1/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2016__A1 _2136_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input87_A gpio_dat_i[21] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2567__A2 _2322_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2801__A _3489_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2520__B _2520_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__D1 _3903_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output243_A _3158_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2947__S _2947_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3632__A _3632_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4339__CLK _4347_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2248__A _2514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3070__C _3600_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _2155_/X _2072_/Y _3470_/X _3314_/X vssd1 vssd1 vccd1 vccd1 _4348_/D sky130_fd_sc_hd__a211o_1
XANTENNA__2682__S _2950_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3079__A _3115_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3861_ _3861_/A _3869_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3862_/A sky130_fd_sc_hd__and3_1
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2812_ _2828_/A _2812_/B _3386_/A vssd1 vssd1 vccd1 vccd1 _2813_/A sky130_fd_sc_hd__and3_2
X_3792_ _3792_/A _3796_/B _3903_/A vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__and3_1
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2743_ _2743_/A vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2558__A2 _3617_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3807__A _3807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2711__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2674_ _3889_/A _4047_/Q _2936_/S vssd1 vssd1 vccd1 vccd1 _3279_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3245__C _3250_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4344_ _4347_/CLK _4344_/D vssd1 vssd1 vccd1 vccd1 _4344_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2191__B1 _2190_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2857__S _2905_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4275_/CLK _4275_/D vssd1 vssd1 vccd1 vccd1 _4275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3691__B1 _4394_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3157_ _3178_/C _4183_/Q _3157_/S vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__mux2_2
XANTENNA__2494__A1 _2406_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2158__A _2158_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2113_/A _2108_/B vssd1 vssd1 vccd1 vccd1 _2346_/A sky130_fd_sc_hd__nand2_4
X_3088_ _3219_/B _4198_/Q _3109_/S vssd1 vssd1 vccd1 vccd1 _3611_/C sky130_fd_sc_hd__mux2_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2039_ _2059_/A vssd1 vssd1 vccd1 vccd1 _2152_/A sky130_fd_sc_hd__buf_2
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3994__B2 _2596_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__A1 _3968_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2549__A2 _2289_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3746__B2 _2396_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3746__A1 _4258_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3717__A _3717_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3452__A _3452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input141_A spi_err_i vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2485__A1 _2283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_13_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A1 _3968_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3985__B2 _2547_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3737__A1 _3765_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4011__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output193_A _3025_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3627__A _3627_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2531__A _2531_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2960__A2 _2133_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3346__B _3346_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4161__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2390_ _4258_/Q vssd1 vssd1 vccd1 vccd1 _2390_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2173__B1 _2172_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3362__A _3362_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4060_ _4326_/CLK _4060_/D vssd1 vssd1 vccd1 vccd1 _4060_/Q sky130_fd_sc_hd__dfxtp_1
X_3011_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__B _3089_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2706__A _2752_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2228__A1 _4285_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1967__D _1967_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3913_ input5/X _3908_/X _3911_/X _3912_/Y vssd1 vssd1 vccd1 vccd1 _4336_/D sky130_fd_sc_hd__a211o_1
X_3844_ _3844_/A vssd1 vssd1 vccd1 vccd1 _4308_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4343__D _4343_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3537__A _3547_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3775_ _3769_/X _3764_/X _3765_/X _2576_/Y _3774_/X vssd1 vssd1 vccd1 vccd1 _4273_/D
+ sky130_fd_sc_hd__o311a_1
X_2726_ _2726_/A _4133_/Q vssd1 vssd1 vccd1 vccd1 _2727_/A sky130_fd_sc_hd__and2_1
XANTENNA__1983__C _2053_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2657_ _3271_/B _4114_/Q _2942_/S vssd1 vssd1 vccd1 vccd1 _3449_/C sky130_fd_sc_hd__mux2_4
X_2588_ _2581_/X _2582_/X _2469_/A _2587_/Y vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3900__A1 _1971_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2164__B1 _4341_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3272__A _3272_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4327_ _4346_/CLK _4327_/D vssd1 vssd1 vccd1 vccd1 _4327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3703__C _3703_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4258_ _4262_/CLK _4258_/D vssd1 vssd1 vccd1 vccd1 _4258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2467__A1 _2465_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ _3209_/A vssd1 vssd1 vccd1 vccd1 _4019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4189_ _4225_/CLK _4189_/D vssd1 vssd1 vccd1 vccd1 _4189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__D _2074_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4034__CLK _4380_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3967__A1 _4365_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4253__D _4253_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3719__A1 _4246_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3719__B2 _3697_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3447__A _3447_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4184__CLK _4262_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3352__C1 _3350_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2155__B1 _4348_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3182__A _3953_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2458__A1 _2262_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2483__A_N _2382_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output206_A _2987_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2526__A _2526_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3121__S _3147_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4163__D _4163_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__A1 _4280_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2630__B2 input95/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__A _3369_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3560_ _3562_/A _3560_/B vssd1 vssd1 vccd1 vccd1 _4175_/D sky130_fd_sc_hd__nor2_1
X_2511_ _2502_/X _2510_/Y _2499_/X _2469_/X vssd1 vssd1 vccd1 vccd1 _2511_/X sky130_fd_sc_hd__o211a_1
X_3491_ _4130_/Q _3488_/X _3489_/X _3490_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _4130_/D
+ sky130_fd_sc_hd__a221o_1
X_2442_ _2380_/X _2438_/Y _2441_/X _2398_/X vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2373_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2373_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2697__A1 _4051_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4112_ _4250_/CLK _4112_/D vssd1 vssd1 vccd1 vccd1 _4112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4043_ _4051_/CLK _4043_/D vssd1 vssd1 vccd1 vccd1 _4043_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4338__D _4338_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3820__A _3820_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4057__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4073__D _4073_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2621__A1 _2427_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2621__B2 _2434_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2082__C1 _1977_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3827_ _3827_/A vssd1 vssd1 vccd1 vccd1 _4301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3758_ _3752_/X _3747_/X _3748_/X _2477_/Y _3757_/X vssd1 vssd1 vccd1 vccd1 _4263_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3267__A _3276_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2171__A _4060_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2709_ _2715_/A _4125_/Q vssd1 vssd1 vccd1 vccd1 _2710_/A sky130_fd_sc_hd__and2_1
X_3689_ _3699_/A _4231_/Q _3703_/C _3689_/D vssd1 vssd1 vccd1 vccd1 _3690_/A sky130_fd_sc_hd__and4_1
Xoutput240 _3075_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[9] sky130_fd_sc_hd__buf_2
Xoutput262 _2736_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput251 _2714_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput284 _2842_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput273 _2685_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput295 _2902_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__3714__B _4243_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3334__C1 _3346_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4248__D _4248_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3730__A _3730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2049__C _3925_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2346__A _2346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input104_A gpio_dat_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__A1 _2581_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2073__C1 _2137_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1966__A3 _1918_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3177__A _3695_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3905__A _3940_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output156_A _2564_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3624__B _3633_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3325__C1 _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3116__S _3144_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3343__C _3343_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3340__A2 _3907_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2143__A3 _3953_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4158__D _4158_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3640__A _3804_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2955__S _2955_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2851__A1 _4096_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2256__A _2452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2991_ _2999_/A _4228_/Q vssd1 vssd1 vccd1 vccd1 _2992_/A sky130_fd_sc_hd__and2_1
XANTENNA__2690__S _2947_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2603__A1 _2581_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ _3953_/A _1942_/B _2023_/A _2022_/A vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__nand4_4
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3087__A _3087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3612_ _3612_/A vssd1 vssd1 vccd1 vccd1 _4198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3543_ _3546_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _4161_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3815__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3474_ _3492_/A _4123_/Q _4002_/B vssd1 vssd1 vccd1 vccd1 _3475_/A sky130_fd_sc_hd__and3_1
XANTENNA__2119__B1 _2517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2425_ _2919_/A _2424_/X _4155_/Q vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__3316__C1 _3315_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3253__C _3253_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2356_ _2356_/A _2356_/B _2356_/C vssd1 vssd1 vccd1 vccd1 _2357_/C sky130_fd_sc_hd__nand3_1
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4068__D _4068_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3550__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2287_ _2529_/A vssd1 vssd1 vccd1 vccd1 _2287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2865__S _2911_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3095__A1 _4200_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _4380_/CLK _4026_/D vssd1 vssd1 vccd1 vccd1 _4026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2070__A2 _3346_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3555__C1 _3547_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2358__B1 _2357_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3725__A _3725_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4222__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3322__A2 _3314_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3460__A _3460_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4372__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2076__A _2076_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2507__C _2507_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2833__A1 _4093_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2804__A _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2597__B1 _2499_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3338__C _3724_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output273_A _2685_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3561__A2 _3447_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3635__A _3635_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3354__B _3774_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__A3 _2272_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2210_ _2210_/A _2210_/B vssd1 vssd1 vccd1 vccd1 _2211_/D sky130_fd_sc_hd__nor2_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2521__B1 _2520_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3190_ _3195_/A _3190_/B _3195_/C _3190_/D vssd1 vssd1 vccd1 vccd1 _3191_/A sky130_fd_sc_hd__or4_1
XFILLER_93_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__A _3383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2141_ _2141_/A vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2072_ input18/X _2072_/B _2078_/C _2078_/D vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2974_ _3326_/D vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2714__A _2714_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2588__B1 _2469_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1925_ _2022_/A _2023_/A vssd1 vssd1 vccd1 vccd1 _1994_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2052__A2 _2015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4351__D _4351_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4245__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3526_ _3526_/A1 _3523_/X _3524_/X _2290_/Y _3562_/A vssd1 vssd1 vccd1 vccd1 _4148_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__2760__A0 _3184_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3457_ _3457_/A _3462_/B _3457_/C vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__or3_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2408_ _2408_/A vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2339_ _2262_/X _2375_/A _2408_/A _2409_/A _2338_/Y vssd1 vssd1 vccd1 vccd1 _2339_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3711__C _3721_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3280__A _3280_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2608__B _2638_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4009_ _4302_/CLK _4009_/D vssd1 vssd1 vccd1 vccd1 _4009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2815__A1 input66/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2291__A2 _2283_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3776__C1 _3772_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3439__B _3459_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4261__D _4261_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2594__A3 _2286_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3455__A _3455_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3174__B _3174_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2074__A_N input20/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A cpu_adr_i[8] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3190__A _3195_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3059__A1 _4190_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4118__CLK _4250_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4268__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4171__D _4171_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2034__A2 _2168_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3782__A2 _3657_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2690_ _3286_/C _4119_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3459_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3365__A _3383_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4360_ _4390_/CLK _4360_/D vssd1 vssd1 vccd1 vccd1 _4360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3311_ _3311_/A vssd1 vssd1 vccd1 vccd1 _4058_/D sky130_fd_sc_hd__clkbuf_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4347_/CLK _4291_/D vssd1 vssd1 vccd1 vccd1 _4291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3242_/A vssd1 vssd1 vccd1 vccd1 _4032_/D sky130_fd_sc_hd__clkbuf_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2709__A _2715_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3173_ _3343_/C vssd1 vssd1 vccd1 vccd1 _3195_/C sky130_fd_sc_hd__clkbuf_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2124_ _4002_/C vssd1 vssd1 vccd1 vccd1 _2579_/A sky130_fd_sc_hd__inv_2
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4346__D _4346_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3250__D _3271_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2055_ _2055_/A _2055_/B vssd1 vssd1 vccd1 vccd1 _2134_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2444__A _2529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3758__C1 _3757_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4081__D _4081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2957_ _4290_/Q input70/X _2957_/S vssd1 vssd1 vccd1 vccd1 _3798_/C sky130_fd_sc_hd__mux2_1
XFILLER_50_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2025__A2 _1970_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2888_ _2888_/A _2901_/B _3418_/C vssd1 vssd1 vccd1 vccd1 _2889_/A sky130_fd_sc_hd__and3_1
XANTENNA__3773__A2 _3767_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2981__A0 _3288_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3275__A _3298_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3509_ _4140_/Q _3308_/A _2767_/A _3490_/A _3504_/X vssd1 vssd1 vccd1 vccd1 _4140_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3930__C1 _3314_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2497__C1 _4372_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4256__D _4256_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2057__C _2057_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1953__B1_N _4337_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2354__A _2514_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3749__C1 _3740_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2016__A2 _2015_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3185__A _3185_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2520__C _2520_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__C1 _3909_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xinput140 spi_dat_i[9] vssd1 vssd1 vccd1 vccd1 _2436_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output236_A _3061_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2529__A _2529_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3124__S _3144_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4166__D _4166_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4090__CLK _4251_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1999__D1 _1965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2264__A _2264_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _3884_/A vssd1 vssd1 vccd1 vccd1 _3879_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2811_ _3208_/C _4089_/Q _2858_/S vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__mux2_2
X_3791_ _3884_/A vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2742_ _2748_/A _4140_/Q vssd1 vssd1 vccd1 vccd1 _2743_/A sky130_fd_sc_hd__and2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2963__B1 _3659_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3807__B _3821_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2711__B _4126_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2673_ _4327_/Q input27/X _2935_/S vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__mux2_4
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3245__D _3245_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4343_ _4347_/CLK _4343_/D vssd1 vssd1 vccd1 vccd1 _4343_/Q sky130_fd_sc_hd__dfxtp_1
X_4274_ _4282_/CLK _4274_/D vssd1 vssd1 vccd1 vccd1 _4274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2191__A1 _2139_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3823__A _3823_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3225_ _3225_/A vssd1 vssd1 vccd1 vccd1 _4026_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2439__A _4260_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2479__C1 _2478_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3691__A1 _4232_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3156_ _2988_/A _2200_/A _3572_/C vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2494__A2 _2407_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2158__B _2158_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3691__B2 _3678_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3087_ _3087_/A vssd1 vssd1 vccd1 vccd1 _3087_/X sky130_fd_sc_hd__clkbuf_1
X_2107_ _2129_/A _2129_/B _4285_/Q vssd1 vssd1 vccd1 vccd1 _2108_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__4076__D _4076_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3979__C1 _3966_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2038_ _2038_/A _2072_/B _2081_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2038_/Y sky130_fd_sc_hd__nand4_2
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3994__A2 _3969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2902__A _2902_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3746__A2 _3734_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2403__C1 _2402_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3989_ _3989_/A _3999_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__and3_1
XANTENNA__3717__B _4245_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2954__A0 _3796_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3131__A0 _3250_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2349__A _2349_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2485__A2 _2483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_input134_A spi_dat_i[3] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__C1 _2246_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3985__A2 _3969_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2084__A _2084_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2812__A _2828_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3737__A2 _3736_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__A _3908_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2945__A0 _4287_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output186_A _3011_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4306__CLK _4371_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3346__C _3346_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2958__S _2958_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3643__A _3643_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2173__A1 input9/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2259__A _2517_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3010_ _3010_/A _4237_/Q vssd1 vssd1 vccd1 vccd1 _3011_/A sky130_fd_sc_hd__and2_1
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__C _3607_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2693__S _2950_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2228__A2 _2130_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2633__C1 _2632_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3912_ _3942_/C _1996_/X _3566_/A vssd1 vssd1 vccd1 vccd1 _3912_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3843_ _3847_/A _3853_/B _3843_/C vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__or3_1
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2722__A _2726_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3818__A _3818_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3774_ _3774_/A vssd1 vssd1 vccd1 vccd1 _3774_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2936__A0 _3874_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2725_ _2725_/A vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1983__D _2081_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2656_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2942_/S sky130_fd_sc_hd__buf_2
XANTENNA__2868__S _2904_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2587_ _2526_/X _2584_/Y _2509_/X _2585_/Y _2586_/Y vssd1 vssd1 vccd1 vccd1 _2587_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__2164__A1 _1952_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3900__A2 _1971_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4326_ _4326_/CLK _4326_/D vssd1 vssd1 vccd1 vccd1 _4326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3703__D _3711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _4284_/CLK _4257_/D vssd1 vssd1 vccd1 vccd1 _4257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4188_ _4284_/CLK _4188_/D vssd1 vssd1 vccd1 vccd1 _4188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3208_ _3221_/A _3227_/B _3208_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3209_/A sky130_fd_sc_hd__and4_1
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3139_ _3151_/A _3142_/B _3646_/C vssd1 vssd1 vccd1 vccd1 _3140_/A sky130_fd_sc_hd__and3_1
XANTENNA__2467__A2 _2411_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3967__A2 _3965_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3719__A2 _3167_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3728__A _3728_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4329__CLK _4346_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2927__A0 _3260_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2560__B1_N _4167_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3447__B _3447_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2778__S _2826_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3463__A _3463_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3352__B1 _3349_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2155__A1 _1971_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__A2 _2452_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__A _2807_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__A2 _2295_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__A _3638_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _3490_/X sky130_fd_sc_hd__clkbuf_2
X_2510_ _2255_/X _2505_/Y _2508_/X _2509_/X vssd1 vssd1 vccd1 vccd1 _2510_/Y sky130_fd_sc_hd__o22ai_4
X_2441_ _2439_/Y _3673_/B _2440_/Y vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3373__A _3373_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2372_ _2579_/A vssd1 vssd1 vccd1 vccd1 _2469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4111_ _4251_/CLK _4111_/D vssd1 vssd1 vccd1 vccd1 _4111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4042_ _4085_/CLK _4042_/D vssd1 vssd1 vccd1 vccd1 _4042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2717__A _2739_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_92_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2606__C1 _4384_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4354__D _4354_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2621__A2 _2428_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2082__B1 _2081_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2452__A _2452_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2909__A0 _4316_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3826_ _3826_/A _3845_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__and3_1
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3757_ _3774_/A vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3267__B _3267_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2708_ _2708_/A vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__clkbuf_1
X_3688_ _4230_/Q _3351_/X _4394_/A _3678_/X _3683_/X vssd1 vssd1 vccd1 vccd1 _4230_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_12_CLK_A clkbuf_2_3_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput252 _2716_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[14] sky130_fd_sc_hd__buf_2
Xoutput230 _3146_/X vssd1 vssd1 vccd1 vccd1 gpio_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput241 _3154_/X vssd1 vssd1 vccd1 vccd1 gpio_sel_o[0] sky130_fd_sc_hd__buf_2
X_2639_ _2637_/Y _2366_/A _2638_/Y vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3334__B1 _3333_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3283__A _3320_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput263 _2738_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput285 _2848_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput274 _2691_/X vssd1 vssd1 vccd1 vccd1 spi_adr_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__3714__C _3721_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xoutput296 _2908_/X vssd1 vssd1 vccd1 vccd1 spi_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__2542__D1 _2541_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4309_ _4371_/CLK _4309_/D vssd1 vssd1 vccd1 vccd1 _4309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_27_CLK_A clkbuf_2_0_0_CLK/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3730__B _3730_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4264__D _4264_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4151__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3458__A _3458_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2612__A2 _2582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2073__B1 _2072_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2362__A _2380_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2081__B _2081_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input62_A cpu_dat_i[5] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3193__A _3193_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3624__C _3624_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3325__B1 _2184_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output149_A _2500_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_94_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output316_A _4395_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4174__D _4174_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _3036_/A vssd1 vssd1 vccd1 vccd1 _2999_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2603__A2 _2582_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3368__A _3368_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2064__B1 _2063_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1941_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1942_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2272__A _2272_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _3611_/A _3611_/B _3611_/C vssd1 vssd1 vccd1 vccd1 _3612_/A sky130_fd_sc_hd__or3_1
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3542_ _2483_/C _3536_/X _3528_/X _2484_/Y _3537_/X vssd1 vssd1 vccd1 vccd1 _4160_/D
+ sky130_fd_sc_hd__a311o_1
X_3473_ _3516_/A vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2119__A1 _2346_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3815__B _3829_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2424_ _2424_/A vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__buf_2
XANTENNA__2119__B2 _2450_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3316__B1 _1947_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2355_ _4180_/Q _2353_/Y _2644_/A _2644_/B vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__a22o_1
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3253__D _3260_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4024__CLK _4085_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4349__D _4349_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3831__A _3831_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3550__B _3550_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2286_ _2286_/A vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__buf_4
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4174__CLK _4177_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4025_ _4051_/CLK _4025_/D vssd1 vssd1 vccd1 vccd1 _4025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4084__D _4084_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2881__S _2905_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3278__A _3293_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2182__A _2182_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3809_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3555__B1 _3524_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2358__A1 _2342_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4259__D _4259_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2357__A _2357_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3491__C1 _3483_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2507__D _2507_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2791__S _2937_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2076__B _2076_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2046__B1 _4065_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2597__A1 _2592_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2092__A _2207_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3188__A _3192_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3338__D _3724_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3916__A _3938_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4047__CLK _4051_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA_output266_A _2745_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3635__B _3635_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3354__C _3376_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4169__D _4169_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2966__S _3335_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A _3651_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2521__A1 _2519_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4197__CLK _4275_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2140_ _2136_/X _3942_/A _4055_/Q vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3370__B _3389_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2267__A _2454_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2071_ _4068_/Q _4070_/Q _2015_/X _2136_/A vssd1 vssd1 vccd1 vccd1 _2076_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2973_ _3343_/C vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2588__A1 _2581_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_1924_ _1924_/A vssd1 vssd1 vccd1 vccd1 _2023_/A sky130_fd_sc_hd__buf_2
XANTENNA__3826__A _3826_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2730__A _2730_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3525_ _3547_/A vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__buf_2
XANTENNA__2760__A1 _4081_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3456_ _3456_/A vssd1 vssd1 vccd1 vccd1 _4117_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4079__D _4079_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2407_ _2407_/A vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2876__S _2886_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3387_ _3387_/A vssd1 vssd1 vccd1 vccd1 _4089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2338_ _2334_/Y _2539_/A _2337_/Y vssd1 vssd1 vccd1 vccd1 _2338_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3711__D _3711_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2269_ _2344_/A vssd1 vssd1 vccd1 vccd1 _2539_/A sky130_fd_sc_hd__buf_4
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2608__C _2638_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_73_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4008_ _4051_/CLK _4008_/D vssd1 vssd1 vccd1 vccd1 _4008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2276__B1 _2275_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2291__A3 _2286_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3776__B1 _3771_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3439__C _3455_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3455__B _3459_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3174__C _3195_/C vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2786__S _2955_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A cpu_adr_i[30] vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2087__A _2087_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3190__B _3190_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2019__B1 _4063_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3646__A _3659_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3519__B1 _3800_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3365__B _3365_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_99_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3310_ _3343_/A _3326_/C _3323_/C _2207_/A vssd1 vssd1 vccd1 vccd1 _3311_/A sky130_fd_sc_hd__or4b_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4290_ _4302_/CLK _4290_/D vssd1 vssd1 vccd1 vccd1 _4290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3241_ _3250_/A _3241_/B _3250_/C _3245_/D vssd1 vssd1 vccd1 vccd1 _3242_/A sky130_fd_sc_hd__or4_1
XANTENNA__3381__A _3381_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2696__S _2953_/S vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_67_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3172_ _3876_/A vssd1 vssd1 vccd1 vccd1 _3195_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2709__B _4125_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2123_ _4391_/Q _2357_/A _3945_/C vssd1 vssd1 vccd1 vccd1 _4002_/C sky130_fd_sc_hd__o21ai_4
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2054_ _1952_/A _2160_/A _4354_/Q vssd1 vssd1 vccd1 vccd1 _3938_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__2725__A _2725_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4212__CLK _4282_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3758__B1 _2477_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4362__D _4362_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2956_ _2704_/A _2133_/A _3361_/A vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2887_ _3241_/B _4102_/Q _2911_/S vssd1 vssd1 vccd1 vccd1 _3418_/C sky130_fd_sc_hd__mux2_1
XANTENNA__2981__A1 _4224_/Q vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3556__A _3558_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__4362__CLK _4390_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3508_ _3508_/A vssd1 vssd1 vccd1 vccd1 _4139_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3930__B1 _3470_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3439_ _3439_/A _3459_/B _3455_/C vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__and3_1
XANTENNA__3291__A _3328_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__2497__B1 _2303_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2057__D _2078_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4272__D _4272_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3749__B1 _2416_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3466__A _3466_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_26_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4074_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2520__D _2520_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__B1 _2028_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2488__B1 _2487_/Y vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput130 spi_dat_i[29] vssd1 vssd1 vccd1 vccd1 _2628_/C sky130_fd_sc_hd__clkbuf_2
Xinput141 spi_err_i vssd1 vssd1 vccd1 vccd1 _2382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output229_A _3143_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4235__CLK _4264_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_64_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1999__C1 _1973_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4182__D _4182_/D vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4385__CLK _4389_/CLK vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _3197_/A vssd1 vssd1 vccd1 vccd1 _2858_/S sky130_fd_sc_hd__buf_2
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _3884_/A sky130_fd_sc_hd__clkbuf_2
X_2741_ _2741_/A vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__clkbuf_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2963__A1 _2197_/X vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_17_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _4280_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2280__A _2418_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3376__A _3376_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XANTENNA__3807__C _3903_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_2672_ _2128_/X _2133_/X _3453_/C vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3912__B1 _3566_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4342_ _4347_/CLK _4342_/D vssd1 vssd1 vccd1 vccd1 _4342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2191__A2 _2864_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_4273_ _4275_/CLK _4273_/D vssd1 vssd1 vccd1 vccd1 _4273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3823__B _3829_/B vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4000__A _4000_/A vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__fakediode_2
X_3224_ _3224_/A _3224_/B _3224_/C _3245_/D vssd1 vssd1 vccd1 vccd1 _3225_/A sky130_fd_sc_hd__or4_1
.ends

