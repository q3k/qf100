magic
tech sky130A
magscale 1 2
timestamp 1647787485
<< viali >>
rect 23673 16609 23707 16643
rect 22937 16541 22971 16575
rect 23397 16541 23431 16575
rect 23489 16541 23523 16575
rect 25145 16541 25179 16575
rect 27537 16541 27571 16575
rect 28549 16541 28583 16575
rect 25412 16473 25446 16507
rect 28273 16473 28307 16507
rect 22753 16405 22787 16439
rect 23673 16405 23707 16439
rect 26525 16405 26559 16439
rect 27353 16405 27387 16439
rect 28371 16405 28405 16439
rect 28457 16405 28491 16439
rect 25605 16201 25639 16235
rect 26341 16133 26375 16167
rect 26985 16133 27019 16167
rect 22385 16065 22419 16099
rect 22652 16065 22686 16099
rect 24225 16065 24259 16099
rect 24481 16065 24515 16099
rect 26065 16065 26099 16099
rect 27169 16065 27203 16099
rect 27261 16065 27295 16099
rect 28273 16065 28307 16099
rect 28529 16065 28563 16099
rect 30461 16065 30495 16099
rect 32137 16065 32171 16099
rect 32321 16065 32355 16099
rect 26341 15997 26375 16031
rect 30205 15997 30239 16031
rect 26157 15929 26191 15963
rect 26985 15929 27019 15963
rect 23765 15861 23799 15895
rect 29653 15861 29687 15895
rect 31585 15861 31619 15895
rect 32137 15861 32171 15895
rect 22845 15657 22879 15691
rect 23029 15657 23063 15691
rect 23489 15657 23523 15691
rect 28917 15657 28951 15691
rect 29929 15657 29963 15691
rect 30757 15657 30791 15691
rect 28825 15589 28859 15623
rect 29009 15521 29043 15555
rect 30849 15521 30883 15555
rect 20637 15453 20671 15487
rect 22477 15453 22511 15487
rect 23489 15453 23523 15487
rect 23765 15453 23799 15487
rect 24593 15453 24627 15487
rect 25053 15453 25087 15487
rect 26893 15453 26927 15487
rect 27160 15453 27194 15487
rect 28733 15453 28767 15487
rect 29929 15453 29963 15487
rect 30113 15453 30147 15487
rect 30573 15453 30607 15487
rect 30665 15453 30699 15487
rect 31309 15453 31343 15487
rect 31576 15453 31610 15487
rect 20904 15385 20938 15419
rect 25298 15385 25332 15419
rect 22017 15317 22051 15351
rect 22845 15317 22879 15351
rect 23673 15317 23707 15351
rect 24409 15317 24443 15351
rect 26433 15317 26467 15351
rect 28273 15317 28307 15351
rect 32689 15317 32723 15351
rect 21833 15113 21867 15147
rect 22753 15113 22787 15147
rect 25605 15113 25639 15147
rect 27813 15113 27847 15147
rect 31401 15113 31435 15147
rect 25421 15045 25455 15079
rect 27629 15045 27663 15079
rect 32137 15045 32171 15079
rect 32337 15045 32371 15079
rect 19892 14977 19926 15011
rect 22017 14977 22051 15011
rect 22937 14977 22971 15011
rect 23121 14977 23155 15011
rect 23213 14977 23247 15011
rect 23857 14977 23891 15011
rect 26249 14977 26283 15011
rect 28457 14977 28491 15011
rect 31125 14977 31159 15011
rect 31217 14977 31251 15011
rect 19625 14909 19659 14943
rect 22293 14909 22327 14943
rect 23673 14909 23707 14943
rect 25053 14909 25087 14943
rect 28273 14909 28307 14943
rect 27261 14841 27295 14875
rect 21005 14773 21039 14807
rect 22201 14773 22235 14807
rect 24041 14773 24075 14807
rect 25421 14773 25455 14807
rect 26065 14773 26099 14807
rect 27629 14773 27663 14807
rect 28641 14773 28675 14807
rect 32321 14773 32355 14807
rect 32505 14773 32539 14807
rect 20545 14569 20579 14603
rect 21925 14569 21959 14603
rect 23397 14569 23431 14603
rect 24777 14569 24811 14603
rect 25421 14569 25455 14603
rect 26709 14569 26743 14603
rect 27353 14569 27387 14603
rect 28641 14569 28675 14603
rect 31125 14569 31159 14603
rect 18429 14501 18463 14535
rect 19717 14433 19751 14467
rect 31217 14433 31251 14467
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 20453 14365 20487 14399
rect 20545 14365 20579 14399
rect 21189 14365 21223 14399
rect 21281 14365 21315 14399
rect 22201 14365 22235 14399
rect 23029 14365 23063 14399
rect 23213 14365 23247 14399
rect 24409 14365 24443 14399
rect 25605 14365 25639 14399
rect 25881 14365 25915 14399
rect 26341 14365 26375 14399
rect 26525 14365 26559 14399
rect 27537 14365 27571 14399
rect 27813 14365 27847 14399
rect 28273 14365 28307 14399
rect 28457 14365 28491 14399
rect 29745 14365 29779 14399
rect 30205 14365 30239 14399
rect 30389 14365 30423 14399
rect 30941 14365 30975 14399
rect 31033 14365 31067 14399
rect 31677 14365 31711 14399
rect 31861 14365 31895 14399
rect 18429 14297 18463 14331
rect 20177 14297 20211 14331
rect 21925 14297 21959 14331
rect 25789 14297 25823 14331
rect 18613 14229 18647 14263
rect 19257 14229 19291 14263
rect 20269 14229 20303 14263
rect 21465 14229 21499 14263
rect 22109 14229 22143 14263
rect 24777 14229 24811 14263
rect 24961 14229 24995 14263
rect 27721 14229 27755 14263
rect 29561 14229 29595 14263
rect 30297 14229 30331 14263
rect 31769 14229 31803 14263
rect 19533 14025 19567 14059
rect 20091 14025 20125 14059
rect 26433 14025 26467 14059
rect 27813 14025 27847 14059
rect 28549 14025 28583 14059
rect 31493 14025 31527 14059
rect 33609 14025 33643 14059
rect 18420 13957 18454 13991
rect 19993 13957 20027 13991
rect 21833 13957 21867 13991
rect 22033 13957 22067 13991
rect 24317 13957 24351 13991
rect 26249 13957 26283 13991
rect 27629 13957 27663 13991
rect 32474 13957 32508 13991
rect 20177 13889 20211 13923
rect 20269 13889 20303 13923
rect 21281 13889 21315 13923
rect 24225 13889 24259 13923
rect 24409 13889 24443 13923
rect 25145 13889 25179 13923
rect 25237 13889 25271 13923
rect 25881 13889 25915 13923
rect 28457 13889 28491 13923
rect 28641 13889 28675 13923
rect 29377 13889 29411 13923
rect 29644 13889 29678 13923
rect 31217 13889 31251 13923
rect 32229 13889 32263 13923
rect 18153 13821 18187 13855
rect 22753 13821 22787 13855
rect 23029 13821 23063 13855
rect 24041 13821 24075 13855
rect 24593 13821 24627 13855
rect 25421 13821 25455 13855
rect 28273 13821 28307 13855
rect 31309 13821 31343 13855
rect 31493 13821 31527 13855
rect 27261 13753 27295 13787
rect 21097 13685 21131 13719
rect 22017 13685 22051 13719
rect 22201 13685 22235 13719
rect 26249 13685 26283 13719
rect 27629 13685 27663 13719
rect 28825 13685 28859 13719
rect 30757 13685 30791 13719
rect 23581 13481 23615 13515
rect 31953 13481 31987 13515
rect 30849 13413 30883 13447
rect 21649 13345 21683 13379
rect 23765 13345 23799 13379
rect 29561 13345 29595 13379
rect 29837 13345 29871 13379
rect 32137 13345 32171 13379
rect 18061 13277 18095 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19717 13277 19751 13311
rect 20913 13277 20947 13311
rect 21189 13277 21223 13311
rect 23489 13277 23523 13311
rect 24869 13277 24903 13311
rect 25145 13277 25179 13311
rect 26433 13277 26467 13311
rect 26525 13277 26559 13311
rect 27537 13277 27571 13311
rect 27804 13277 27838 13311
rect 31033 13277 31067 13311
rect 31861 13277 31895 13311
rect 21916 13209 21950 13243
rect 26157 13209 26191 13243
rect 31125 13209 31159 13243
rect 17877 13141 17911 13175
rect 18613 13141 18647 13175
rect 19809 13141 19843 13175
rect 20729 13141 20763 13175
rect 21097 13141 21131 13175
rect 23029 13141 23063 13175
rect 23765 13141 23799 13175
rect 26341 13141 26375 13175
rect 26709 13141 26743 13175
rect 28917 13141 28951 13175
rect 31217 13141 31251 13175
rect 31401 13141 31435 13175
rect 32137 13141 32171 13175
rect 22201 12937 22235 12971
rect 22385 12937 22419 12971
rect 24685 12937 24719 12971
rect 25145 12937 25179 12971
rect 25881 12937 25915 12971
rect 28641 12937 28675 12971
rect 30941 12937 30975 12971
rect 32505 12937 32539 12971
rect 19257 12869 19291 12903
rect 23572 12869 23606 12903
rect 30573 12869 30607 12903
rect 30789 12869 30823 12903
rect 9697 12801 9731 12835
rect 10517 12801 10551 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 18153 12801 18187 12835
rect 19901 12801 19935 12835
rect 23305 12801 23339 12835
rect 25329 12801 25363 12835
rect 26157 12801 26191 12835
rect 26249 12801 26283 12835
rect 27353 12801 27387 12835
rect 28825 12801 28859 12835
rect 29009 12801 29043 12835
rect 29837 12801 29871 12835
rect 29929 12801 29963 12835
rect 31401 12801 31435 12835
rect 31585 12801 31619 12835
rect 32321 12801 32355 12835
rect 32413 12801 32447 12835
rect 33793 12801 33827 12835
rect 18429 12733 18463 12767
rect 18889 12733 18923 12767
rect 20177 12733 20211 12767
rect 21833 12733 21867 12767
rect 26065 12733 26099 12767
rect 26341 12733 26375 12767
rect 27629 12733 27663 12767
rect 28917 12733 28951 12767
rect 29101 12733 29135 12767
rect 33609 12733 33643 12767
rect 33701 12733 33735 12767
rect 33885 12733 33919 12767
rect 18337 12665 18371 12699
rect 32137 12665 32171 12699
rect 9505 12597 9539 12631
rect 10333 12597 10367 12631
rect 17417 12597 17451 12631
rect 18245 12597 18279 12631
rect 19257 12597 19291 12631
rect 19441 12597 19475 12631
rect 22201 12597 22235 12631
rect 30113 12597 30147 12631
rect 30757 12597 30791 12631
rect 31401 12597 31435 12631
rect 32689 12597 32723 12631
rect 33425 12597 33459 12631
rect 9965 12393 9999 12427
rect 16405 12393 16439 12427
rect 19901 12393 19935 12427
rect 24409 12393 24443 12427
rect 28733 12393 28767 12427
rect 30021 12393 30055 12427
rect 18337 12325 18371 12359
rect 19349 12325 19383 12359
rect 27445 12325 27479 12359
rect 6745 12257 6779 12291
rect 9597 12257 9631 12291
rect 23305 12257 23339 12291
rect 24593 12257 24627 12291
rect 24777 12257 24811 12291
rect 30113 12257 30147 12291
rect 6929 12189 6963 12223
rect 7849 12189 7883 12223
rect 9137 12189 9171 12223
rect 9781 12189 9815 12223
rect 11345 12189 11379 12223
rect 12081 12189 12115 12223
rect 14565 12189 14599 12223
rect 16221 12189 16255 12223
rect 16957 12189 16991 12223
rect 17224 12189 17258 12223
rect 19625 12189 19659 12223
rect 20637 12189 20671 12223
rect 23029 12189 23063 12223
rect 24685 12189 24719 12223
rect 24869 12189 24903 12223
rect 25605 12189 25639 12223
rect 27721 12189 27755 12223
rect 29837 12189 29871 12223
rect 29929 12189 29963 12223
rect 30757 12189 30791 12223
rect 31217 12189 31251 12223
rect 33057 12189 33091 12223
rect 33333 12189 33367 12223
rect 10517 12121 10551 12155
rect 14749 12121 14783 12155
rect 20904 12121 20938 12155
rect 25872 12121 25906 12155
rect 27445 12121 27479 12155
rect 28641 12121 28675 12155
rect 31484 12121 31518 12155
rect 7113 12053 7147 12087
rect 7665 12053 7699 12087
rect 8953 12053 8987 12087
rect 10609 12053 10643 12087
rect 11161 12053 11195 12087
rect 11897 12053 11931 12087
rect 19533 12053 19567 12087
rect 19717 12053 19751 12087
rect 22017 12053 22051 12087
rect 26985 12053 27019 12087
rect 27629 12053 27663 12087
rect 30573 12053 30607 12087
rect 32597 12053 32631 12087
rect 8585 11849 8619 11883
rect 22109 11849 22143 11883
rect 22385 11849 22419 11883
rect 22937 11849 22971 11883
rect 30205 11849 30239 11883
rect 31033 11849 31067 11883
rect 11774 11781 11808 11815
rect 16037 11781 16071 11815
rect 17202 11781 17236 11815
rect 29092 11781 29126 11815
rect 5825 11713 5859 11747
rect 6377 11713 6411 11747
rect 6633 11713 6667 11747
rect 8401 11713 8435 11747
rect 9137 11713 9171 11747
rect 9393 11713 9427 11747
rect 11529 11713 11563 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 14657 11713 14691 11747
rect 14841 11713 14875 11747
rect 15485 11713 15519 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 19349 11713 19383 11747
rect 19616 11713 19650 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 23673 11713 23707 11747
rect 24409 11713 24443 11747
rect 24676 11713 24710 11747
rect 26433 11713 26467 11747
rect 26985 11713 27019 11747
rect 27241 11713 27275 11747
rect 28825 11713 28859 11747
rect 30849 11713 30883 11747
rect 32321 11713 32355 11747
rect 33057 11713 33091 11747
rect 33313 11713 33347 11747
rect 34897 11713 34931 11747
rect 35153 11713 35187 11747
rect 8217 11645 8251 11679
rect 14105 11645 14139 11679
rect 16957 11645 16991 11679
rect 30665 11645 30699 11679
rect 32597 11645 32631 11679
rect 5641 11577 5675 11611
rect 21833 11577 21867 11611
rect 32137 11577 32171 11611
rect 7757 11509 7791 11543
rect 10517 11509 10551 11543
rect 12909 11509 12943 11543
rect 13369 11509 13403 11543
rect 14749 11509 14783 11543
rect 15301 11509 15335 11543
rect 18337 11509 18371 11543
rect 20729 11509 20763 11543
rect 23489 11509 23523 11543
rect 25789 11509 25823 11543
rect 26249 11509 26283 11543
rect 28365 11509 28399 11543
rect 32505 11509 32539 11543
rect 34437 11509 34471 11543
rect 36277 11509 36311 11543
rect 8401 11305 8435 11339
rect 12449 11305 12483 11339
rect 14473 11305 14507 11339
rect 18061 11305 18095 11339
rect 20545 11305 20579 11339
rect 22753 11305 22787 11339
rect 24685 11305 24719 11339
rect 25053 11305 25087 11339
rect 26985 11305 27019 11339
rect 27353 11305 27387 11339
rect 29929 11305 29963 11339
rect 30113 11305 30147 11339
rect 33977 11305 34011 11339
rect 17325 11237 17359 11271
rect 26341 11237 26375 11271
rect 7021 11169 7055 11203
rect 9137 11169 9171 11203
rect 10425 11169 10459 11203
rect 18429 11169 18463 11203
rect 25677 11169 25711 11203
rect 27445 11169 27479 11203
rect 29561 11169 29595 11203
rect 30941 11169 30975 11203
rect 32689 11169 32723 11203
rect 5181 11101 5215 11135
rect 7288 11101 7322 11135
rect 9413 11101 9447 11135
rect 12265 11101 12299 11135
rect 14105 11101 14139 11135
rect 14381 11101 14415 11135
rect 15117 11101 15151 11135
rect 15384 11101 15418 11135
rect 17601 11101 17635 11135
rect 18245 11101 18279 11135
rect 18337 11101 18371 11135
rect 18521 11101 18555 11135
rect 19257 11101 19291 11135
rect 19533 11101 19567 11135
rect 20729 11101 20763 11135
rect 21189 11101 21223 11135
rect 21373 11101 21407 11135
rect 23397 11101 23431 11135
rect 24869 11101 24903 11135
rect 25145 11101 25179 11135
rect 25881 11101 25915 11135
rect 26525 11101 26559 11135
rect 27169 11101 27203 11135
rect 28089 11101 28123 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 30757 11101 30791 11135
rect 31033 11101 31067 11135
rect 31769 11101 31803 11135
rect 32965 11101 32999 11135
rect 33977 11101 34011 11135
rect 34161 11101 34195 11135
rect 5448 11033 5482 11067
rect 10692 11033 10726 11067
rect 13369 11033 13403 11067
rect 13553 11033 13587 11067
rect 17325 11033 17359 11067
rect 21281 11033 21315 11067
rect 22385 11033 22419 11067
rect 22569 11033 22603 11067
rect 23581 11033 23615 11067
rect 23765 11033 23799 11067
rect 25605 11033 25639 11067
rect 28549 11033 28583 11067
rect 29929 11033 29963 11067
rect 31585 11033 31619 11067
rect 6561 10965 6595 10999
rect 11805 10965 11839 10999
rect 14657 10965 14691 10999
rect 16497 10965 16531 10999
rect 17509 10965 17543 10999
rect 25789 10965 25823 10999
rect 27905 10965 27939 10999
rect 28917 10965 28951 10999
rect 30573 10965 30607 10999
rect 5641 10761 5675 10795
rect 7297 10761 7331 10795
rect 9965 10761 9999 10795
rect 10977 10761 11011 10795
rect 13737 10761 13771 10795
rect 17693 10761 17727 10795
rect 18981 10761 19015 10795
rect 25697 10761 25731 10795
rect 30941 10761 30975 10795
rect 32965 10761 32999 10795
rect 33701 10761 33735 10795
rect 8125 10693 8159 10727
rect 11713 10693 11747 10727
rect 11897 10693 11931 10727
rect 12602 10693 12636 10727
rect 17509 10693 17543 10727
rect 18337 10693 18371 10727
rect 22661 10693 22695 10727
rect 22753 10693 22787 10727
rect 29828 10693 29862 10727
rect 5825 10625 5859 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 7113 10625 7147 10659
rect 7941 10625 7975 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 9781 10625 9815 10659
rect 10609 10625 10643 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 12357 10625 12391 10659
rect 14197 10625 14231 10659
rect 15485 10625 15519 10659
rect 15761 10625 15795 10659
rect 16681 10625 16715 10659
rect 16865 10625 16899 10659
rect 17785 10625 17819 10659
rect 19257 10625 19291 10659
rect 19349 10625 19383 10659
rect 19441 10625 19475 10659
rect 21189 10625 21223 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22477 10625 22511 10659
rect 22845 10625 22879 10659
rect 23673 10625 23707 10659
rect 23857 10625 23891 10659
rect 24869 10625 24903 10659
rect 25605 10625 25639 10659
rect 26249 10625 26283 10659
rect 26433 10625 26467 10659
rect 27077 10625 27111 10659
rect 28181 10625 28215 10659
rect 28917 10625 28951 10659
rect 29561 10625 29595 10659
rect 31585 10625 31619 10659
rect 32321 10625 32355 10659
rect 32781 10625 32815 10659
rect 33057 10625 33091 10659
rect 33517 10625 33551 10659
rect 33793 10625 33827 10659
rect 34253 10625 34287 10659
rect 34529 10625 34563 10659
rect 35725 10625 35759 10659
rect 7757 10557 7791 10591
rect 9597 10557 9631 10591
rect 14473 10557 14507 10591
rect 15945 10557 15979 10591
rect 16129 10557 16163 10591
rect 19165 10557 19199 10591
rect 19993 10557 20027 10591
rect 23949 10557 23983 10591
rect 9137 10489 9171 10523
rect 17509 10489 17543 10523
rect 18521 10489 18555 10523
rect 20361 10489 20395 10523
rect 21005 10489 21039 10523
rect 26249 10489 26283 10523
rect 29101 10489 29135 10523
rect 32781 10489 32815 10523
rect 33517 10489 33551 10523
rect 16773 10421 16807 10455
rect 20453 10421 20487 10455
rect 21833 10421 21867 10455
rect 23029 10421 23063 10455
rect 23489 10421 23523 10455
rect 24961 10421 24995 10455
rect 27169 10421 27203 10455
rect 28273 10421 28307 10455
rect 31401 10421 31435 10455
rect 32137 10421 32171 10455
rect 35541 10421 35575 10455
rect 7113 10217 7147 10251
rect 8217 10217 8251 10251
rect 9505 10217 9539 10251
rect 11253 10217 11287 10251
rect 13369 10217 13403 10251
rect 15761 10217 15795 10251
rect 16865 10217 16899 10251
rect 17601 10217 17635 10251
rect 22937 10217 22971 10251
rect 29929 10217 29963 10251
rect 36001 10217 36035 10251
rect 10333 10149 10367 10183
rect 18337 10149 18371 10183
rect 21649 10149 21683 10183
rect 25881 10149 25915 10183
rect 28457 10149 28491 10183
rect 30941 10149 30975 10183
rect 26617 10081 26651 10115
rect 31401 10081 31435 10115
rect 33517 10081 33551 10115
rect 5273 10013 5307 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7665 10013 7699 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 8953 10013 8987 10047
rect 9321 10013 9355 10047
rect 10977 10013 11011 10047
rect 11069 10013 11103 10047
rect 11345 10013 11379 10047
rect 11897 10013 11931 10047
rect 13277 10013 13311 10047
rect 14473 10013 14507 10047
rect 14657 10013 14691 10047
rect 14841 10013 14875 10047
rect 15393 10013 15427 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16497 10013 16531 10047
rect 16681 10013 16715 10047
rect 18153 10013 18187 10047
rect 20361 10013 20395 10047
rect 22569 10013 22603 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 23857 10013 23891 10047
rect 24409 10013 24443 10047
rect 24557 10013 24591 10047
rect 24685 10013 24719 10047
rect 24915 10013 24949 10047
rect 25789 10013 25823 10047
rect 25973 10013 26007 10047
rect 26884 10013 26918 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 30205 10013 30239 10047
rect 30757 10013 30791 10047
rect 31585 10013 31619 10047
rect 31769 10013 31803 10047
rect 32413 10013 32447 10047
rect 33057 10013 33091 10047
rect 33149 10013 33183 10047
rect 33977 10013 34011 10047
rect 34161 10013 34195 10047
rect 35173 10013 35207 10047
rect 35909 10013 35943 10047
rect 5457 9945 5491 9979
rect 6745 9945 6779 9979
rect 7849 9945 7883 9979
rect 9137 9945 9171 9979
rect 9229 9945 9263 9979
rect 10149 9945 10183 9979
rect 14289 9945 14323 9979
rect 17509 9945 17543 9979
rect 19717 9945 19751 9979
rect 22753 9945 22787 9979
rect 24777 9945 24811 9979
rect 29929 9945 29963 9979
rect 32873 9945 32907 9979
rect 5641 9877 5675 9911
rect 10793 9877 10827 9911
rect 12081 9877 12115 9911
rect 14565 9877 14599 9911
rect 15577 9877 15611 9911
rect 19809 9877 19843 9911
rect 25053 9877 25087 9911
rect 27997 9877 28031 9911
rect 30113 9877 30147 9911
rect 32229 9877 32263 9911
rect 33333 9877 33367 9911
rect 33425 9877 33459 9911
rect 34069 9877 34103 9911
rect 35265 9877 35299 9911
rect 17233 9673 17267 9707
rect 25421 9673 25455 9707
rect 34529 9673 34563 9707
rect 15669 9605 15703 9639
rect 18236 9605 18270 9639
rect 24308 9605 24342 9639
rect 26249 9605 26283 9639
rect 30021 9605 30055 9639
rect 32382 9605 32416 9639
rect 4445 9537 4479 9571
rect 4712 9537 4746 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6653 9537 6687 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 8677 9537 8711 9571
rect 9781 9537 9815 9571
rect 10793 9537 10827 9571
rect 11621 9537 11655 9571
rect 13001 9537 13035 9571
rect 13369 9537 13403 9571
rect 13737 9537 13771 9571
rect 14381 9537 14415 9571
rect 14657 9537 14691 9571
rect 15945 9537 15979 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17095 9537 17129 9571
rect 20361 9537 20395 9571
rect 20545 9537 20579 9571
rect 21005 9537 21039 9571
rect 22201 9537 22235 9571
rect 22468 9537 22502 9571
rect 24041 9537 24075 9571
rect 25881 9537 25915 9571
rect 26065 9537 26099 9571
rect 26985 9537 27019 9571
rect 27169 9537 27203 9571
rect 27988 9537 28022 9571
rect 30205 9537 30239 9571
rect 30757 9537 30791 9571
rect 31401 9537 31435 9571
rect 31585 9537 31619 9571
rect 34253 9537 34287 9571
rect 34391 9537 34425 9571
rect 35081 9537 35115 9571
rect 35265 9537 35299 9571
rect 35357 9537 35391 9571
rect 35817 9537 35851 9571
rect 36001 9537 36035 9571
rect 8769 9469 8803 9503
rect 9505 9469 9539 9503
rect 11897 9469 11931 9503
rect 15761 9469 15795 9503
rect 17969 9469 18003 9503
rect 27721 9469 27755 9503
rect 32137 9469 32171 9503
rect 34161 9469 34195 9503
rect 34621 9469 34655 9503
rect 6837 9401 6871 9435
rect 8217 9401 8251 9435
rect 13185 9401 13219 9435
rect 21097 9401 21131 9435
rect 5825 9333 5859 9367
rect 6377 9333 6411 9367
rect 8677 9333 8711 9367
rect 9045 9333 9079 9367
rect 10885 9333 10919 9367
rect 15761 9333 15795 9367
rect 16129 9333 16163 9367
rect 19349 9333 19383 9367
rect 23581 9333 23615 9367
rect 26985 9333 27019 9367
rect 29101 9333 29135 9367
rect 30849 9333 30883 9367
rect 31401 9333 31435 9367
rect 33517 9333 33551 9367
rect 33977 9333 34011 9367
rect 35173 9333 35207 9367
rect 35817 9333 35851 9367
rect 5733 9129 5767 9163
rect 6193 9129 6227 9163
rect 8033 9129 8067 9163
rect 8401 9129 8435 9163
rect 10609 9129 10643 9163
rect 11989 9129 12023 9163
rect 13553 9129 13587 9163
rect 14105 9129 14139 9163
rect 14473 9129 14507 9163
rect 16037 9129 16071 9163
rect 19901 9129 19935 9163
rect 23673 9129 23707 9163
rect 32045 9129 32079 9163
rect 32229 9129 32263 9163
rect 33977 9129 34011 9163
rect 34161 9129 34195 9163
rect 28733 9061 28767 9095
rect 6653 8993 6687 9027
rect 8033 8993 8067 9027
rect 9505 8993 9539 9027
rect 11069 8993 11103 9027
rect 15189 8993 15223 9027
rect 22293 8993 22327 9027
rect 24961 8993 24995 9027
rect 26801 8993 26835 9027
rect 29653 8993 29687 9027
rect 4353 8925 4387 8959
rect 6377 8925 6411 8959
rect 6469 8925 6503 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 8217 8925 8251 8959
rect 9229 8925 9263 8959
rect 10793 8925 10827 8959
rect 10885 8925 10919 8959
rect 11161 8925 11195 8959
rect 11621 8925 11655 8959
rect 11805 8925 11839 8959
rect 12449 8925 12483 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 15393 8925 15427 8959
rect 15945 8925 15979 8959
rect 16681 8925 16715 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 20131 8925 20165 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 25228 8925 25262 8959
rect 27077 8925 27111 8959
rect 28089 8925 28123 8959
rect 28237 8925 28271 8959
rect 28457 8925 28491 8959
rect 28554 8925 28588 8959
rect 29920 8925 29954 8959
rect 32873 8925 32907 8959
rect 32965 8925 32999 8959
rect 33333 8925 33367 8959
rect 34713 8925 34747 8959
rect 4620 8857 4654 8891
rect 7941 8857 7975 8891
rect 13185 8857 13219 8891
rect 13369 8857 13403 8891
rect 15117 8857 15151 8891
rect 16926 8857 16960 8891
rect 18613 8857 18647 8891
rect 22560 8857 22594 8891
rect 28365 8857 28399 8891
rect 31861 8857 31895 8891
rect 33793 8857 33827 8891
rect 33993 8857 34027 8891
rect 34958 8857 34992 8891
rect 7205 8789 7239 8823
rect 12633 8789 12667 8823
rect 15301 8789 15335 8823
rect 18061 8789 18095 8823
rect 19349 8789 19383 8823
rect 21005 8789 21039 8823
rect 26341 8789 26375 8823
rect 31033 8789 31067 8823
rect 32071 8789 32105 8823
rect 32689 8789 32723 8823
rect 33149 8789 33183 8823
rect 33241 8789 33275 8823
rect 36093 8789 36127 8823
rect 4629 8585 4663 8619
rect 6377 8585 6411 8619
rect 8953 8585 8987 8619
rect 21189 8585 21223 8619
rect 24133 8585 24167 8619
rect 30481 8585 30515 8619
rect 34259 8585 34293 8619
rect 14657 8517 14691 8551
rect 19502 8517 19536 8551
rect 22017 8517 22051 8551
rect 25973 8517 26007 8551
rect 29029 8517 29063 8551
rect 32229 8517 32263 8551
rect 34161 8517 34195 8551
rect 34345 8517 34379 8551
rect 34989 8517 35023 8551
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 7573 8449 7607 8483
rect 7840 8449 7874 8483
rect 9413 8449 9447 8483
rect 9597 8449 9631 8483
rect 10425 8449 10459 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 12541 8449 12575 8483
rect 13369 8449 13403 8483
rect 14473 8449 14507 8483
rect 15301 8449 15335 8483
rect 15577 8449 15611 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 17693 8449 17727 8483
rect 18797 8449 18831 8483
rect 21097 8449 21131 8483
rect 21833 8449 21867 8483
rect 22101 8449 22135 8483
rect 22201 8449 22235 8483
rect 23029 8449 23063 8483
rect 23489 8449 23523 8483
rect 23582 8449 23616 8483
rect 23765 8449 23799 8483
rect 23857 8449 23891 8483
rect 23995 8449 24029 8483
rect 24685 8449 24719 8483
rect 25605 8449 25639 8483
rect 25753 8449 25787 8483
rect 25881 8449 25915 8483
rect 26111 8449 26145 8483
rect 27537 8449 27571 8483
rect 27685 8449 27719 8483
rect 27813 8449 27847 8483
rect 27905 8449 27939 8483
rect 28043 8449 28077 8483
rect 28630 8449 28664 8483
rect 28789 8449 28823 8483
rect 28917 8449 28951 8483
rect 29106 8449 29140 8483
rect 30478 8449 30512 8483
rect 30849 8449 30883 8483
rect 31401 8449 31435 8483
rect 31585 8449 31619 8483
rect 33333 8449 33367 8483
rect 34437 8449 34471 8483
rect 34897 8449 34931 8483
rect 35725 8449 35759 8483
rect 15393 8381 15427 8415
rect 17233 8381 17267 8415
rect 19257 8381 19291 8415
rect 30941 8381 30975 8415
rect 32689 8381 32723 8415
rect 33425 8381 33459 8415
rect 33517 8381 33551 8415
rect 33609 8381 33643 8415
rect 5733 8313 5767 8347
rect 9781 8313 9815 8347
rect 14841 8313 14875 8347
rect 15761 8313 15795 8347
rect 18061 8313 18095 8347
rect 18153 8313 18187 8347
rect 20637 8313 20671 8347
rect 22385 8313 22419 8347
rect 22845 8313 22879 8347
rect 24869 8313 24903 8347
rect 26249 8313 26283 8347
rect 28181 8313 28215 8347
rect 29285 8313 29319 8347
rect 31401 8313 31435 8347
rect 32597 8313 32631 8347
rect 33149 8313 33183 8347
rect 5273 8245 5307 8279
rect 10517 8245 10551 8279
rect 12725 8245 12759 8279
rect 13461 8245 13495 8279
rect 15577 8245 15611 8279
rect 16773 8245 16807 8279
rect 18613 8245 18647 8279
rect 30297 8245 30331 8279
rect 35541 8245 35575 8279
rect 5549 8041 5583 8075
rect 8033 8041 8067 8075
rect 13369 8041 13403 8075
rect 17325 8041 17359 8075
rect 17969 8041 18003 8075
rect 18245 8041 18279 8075
rect 19349 8041 19383 8075
rect 23857 8041 23891 8075
rect 24593 8041 24627 8075
rect 25881 8041 25915 8075
rect 26525 8041 26559 8075
rect 28457 8041 28491 8075
rect 30021 7973 30055 8007
rect 6653 7905 6687 7939
rect 9229 7905 9263 7939
rect 27261 7905 27295 7939
rect 28089 7905 28123 7939
rect 32321 7905 32355 7939
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 6193 7837 6227 7871
rect 11345 7837 11379 7871
rect 14105 7837 14139 7871
rect 15945 7837 15979 7871
rect 17785 7837 17819 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 20085 7837 20119 7871
rect 21005 7837 21039 7871
rect 21189 7837 21223 7871
rect 22477 7837 22511 7871
rect 24409 7837 24443 7871
rect 25513 7837 25547 7871
rect 25697 7837 25731 7871
rect 27445 7837 27479 7871
rect 28273 7837 28307 7871
rect 29837 7837 29871 7871
rect 30573 7837 30607 7871
rect 30665 7837 30699 7871
rect 30941 7837 30975 7871
rect 31125 7837 31159 7871
rect 32045 7837 32079 7871
rect 32137 7837 32171 7871
rect 32413 7837 32447 7871
rect 33793 7837 33827 7871
rect 34897 7837 34931 7871
rect 35357 7837 35391 7871
rect 35541 7837 35575 7871
rect 36185 7837 36219 7871
rect 6920 7769 6954 7803
rect 9474 7769 9508 7803
rect 11612 7769 11646 7803
rect 13277 7769 13311 7803
rect 14372 7769 14406 7803
rect 16212 7769 16246 7803
rect 21649 7769 21683 7803
rect 21833 7769 21867 7803
rect 22722 7769 22756 7803
rect 26433 7769 26467 7803
rect 30849 7769 30883 7803
rect 32965 7769 32999 7803
rect 35449 7769 35483 7803
rect 6009 7701 6043 7735
rect 10609 7701 10643 7735
rect 12725 7701 12759 7735
rect 15485 7701 15519 7735
rect 20269 7701 20303 7735
rect 21189 7701 21223 7735
rect 22017 7701 22051 7735
rect 27629 7701 27663 7735
rect 31861 7701 31895 7735
rect 33057 7701 33091 7735
rect 33609 7701 33643 7735
rect 34713 7701 34747 7735
rect 36001 7701 36035 7735
rect 9137 7497 9171 7531
rect 13553 7497 13587 7531
rect 15025 7497 15059 7531
rect 18245 7497 18279 7531
rect 21097 7497 21131 7531
rect 28457 7497 28491 7531
rect 29101 7497 29135 7531
rect 31217 7497 31251 7531
rect 5457 7429 5491 7463
rect 6561 7429 6595 7463
rect 8769 7429 8803 7463
rect 12081 7429 12115 7463
rect 13185 7429 13219 7463
rect 14013 7429 14047 7463
rect 17110 7429 17144 7463
rect 23305 7429 23339 7463
rect 26249 7429 26283 7463
rect 34980 7429 35014 7463
rect 5641 7361 5675 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 8125 7361 8159 7395
rect 8585 7361 8619 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9873 7361 9907 7395
rect 10057 7361 10091 7395
rect 10149 7361 10183 7395
rect 10241 7361 10275 7395
rect 12265 7361 12299 7395
rect 13369 7361 13403 7395
rect 14197 7361 14231 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 15210 7361 15244 7395
rect 15301 7361 15335 7395
rect 15577 7361 15611 7395
rect 16865 7361 16899 7395
rect 19073 7361 19107 7395
rect 19257 7361 19291 7395
rect 19625 7361 19659 7395
rect 20269 7361 20303 7395
rect 20453 7361 20487 7395
rect 21281 7361 21315 7395
rect 21833 7361 21867 7395
rect 22293 7361 22327 7395
rect 22661 7361 22695 7395
rect 22845 7361 22879 7395
rect 23489 7361 23523 7395
rect 23581 7361 23615 7395
rect 25053 7361 25087 7395
rect 25421 7361 25455 7395
rect 25605 7361 25639 7395
rect 27344 7361 27378 7395
rect 28917 7361 28951 7395
rect 29837 7361 29871 7395
rect 30104 7361 30138 7395
rect 32597 7361 32631 7395
rect 32864 7361 32898 7395
rect 34713 7361 34747 7395
rect 18797 7293 18831 7327
rect 19533 7293 19567 7327
rect 22109 7293 22143 7327
rect 24593 7293 24627 7327
rect 25145 7293 25179 7327
rect 27077 7293 27111 7327
rect 7021 7225 7055 7259
rect 8033 7225 8067 7259
rect 12449 7225 12483 7259
rect 18889 7225 18923 7259
rect 21925 7225 21959 7259
rect 24685 7225 24719 7259
rect 26433 7225 26467 7259
rect 5825 7157 5859 7191
rect 7573 7157 7607 7191
rect 10425 7157 10459 7191
rect 14473 7157 14507 7191
rect 15485 7157 15519 7191
rect 20269 7157 20303 7191
rect 23305 7157 23339 7191
rect 33977 7157 34011 7191
rect 36093 7157 36127 7191
rect 6653 6953 6687 6987
rect 21925 6953 21959 6987
rect 22937 6953 22971 6987
rect 23489 6953 23523 6987
rect 26801 6953 26835 6987
rect 33057 6953 33091 6987
rect 35909 6953 35943 6987
rect 16221 6885 16255 6919
rect 16773 6885 16807 6919
rect 24501 6885 24535 6919
rect 30021 6885 30055 6919
rect 5273 6817 5307 6851
rect 7481 6817 7515 6851
rect 9321 6817 9355 6851
rect 9781 6817 9815 6851
rect 11345 6817 11379 6851
rect 12633 6817 12667 6851
rect 13093 6817 13127 6851
rect 15393 6817 15427 6851
rect 18061 6817 18095 6851
rect 20545 6817 20579 6851
rect 23029 6817 23063 6851
rect 24409 6817 24443 6851
rect 24777 6817 24811 6851
rect 31217 6817 31251 6851
rect 31677 6817 31711 6851
rect 7113 6749 7147 6783
rect 8309 6749 8343 6783
rect 9045 6749 9079 6783
rect 9137 6749 9171 6783
rect 10057 6749 10091 6783
rect 11621 6749 11655 6783
rect 12817 6749 12851 6783
rect 12969 6749 13003 6783
rect 13185 6749 13219 6783
rect 14565 6749 14599 6783
rect 15025 6749 15059 6783
rect 16037 6749 16071 6783
rect 16681 6749 16715 6783
rect 16865 6749 16899 6783
rect 17969 6749 18003 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 22510 6749 22544 6783
rect 23489 6749 23523 6783
rect 23673 6749 23707 6783
rect 24869 6749 24903 6783
rect 25237 6749 25271 6783
rect 25421 6749 25455 6783
rect 26341 6749 26375 6783
rect 26801 6749 26835 6783
rect 26985 6749 27019 6783
rect 27813 6749 27847 6783
rect 28457 6749 28491 6783
rect 29745 6749 29779 6783
rect 29929 6749 29963 6783
rect 30205 6749 30239 6783
rect 30481 6749 30515 6783
rect 31944 6749 31978 6783
rect 33701 6749 33735 6783
rect 34897 6749 34931 6783
rect 35265 6749 35299 6783
rect 36093 6725 36127 6759
rect 36737 6749 36771 6783
rect 37381 6749 37415 6783
rect 5540 6681 5574 6715
rect 7297 6681 7331 6715
rect 14381 6681 14415 6715
rect 15209 6681 15243 6715
rect 18245 6681 18279 6715
rect 18337 6681 18371 6715
rect 20812 6681 20846 6715
rect 27629 6681 27663 6715
rect 27997 6681 28031 6715
rect 31033 6681 31067 6715
rect 35081 6681 35115 6715
rect 35173 6681 35207 6715
rect 8125 6613 8159 6647
rect 19257 6613 19291 6647
rect 19901 6613 19935 6647
rect 22385 6613 22419 6647
rect 22569 6613 22603 6647
rect 26157 6613 26191 6647
rect 28641 6613 28675 6647
rect 33517 6613 33551 6647
rect 35449 6613 35483 6647
rect 36553 6613 36587 6647
rect 37197 6613 37231 6647
rect 4353 6409 4387 6443
rect 4997 6409 5031 6443
rect 6377 6409 6411 6443
rect 16037 6409 16071 6443
rect 17141 6409 17175 6443
rect 19809 6409 19843 6443
rect 30481 6409 30515 6443
rect 34713 6409 34747 6443
rect 35725 6409 35759 6443
rect 36553 6409 36587 6443
rect 8953 6341 8987 6375
rect 12081 6341 12115 6375
rect 15945 6341 15979 6375
rect 18696 6341 18730 6375
rect 22845 6341 22879 6375
rect 27261 6341 27295 6375
rect 32321 6341 32355 6375
rect 34345 6341 34379 6375
rect 35357 6341 35391 6375
rect 35449 6341 35483 6375
rect 36185 6341 36219 6375
rect 4537 6273 4571 6307
rect 5181 6273 5215 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 7573 6273 7607 6307
rect 8217 6273 8251 6307
rect 9597 6273 9631 6307
rect 11897 6273 11931 6307
rect 12992 6273 13026 6307
rect 14565 6273 14599 6307
rect 14749 6273 14783 6307
rect 16681 6273 16715 6307
rect 17785 6273 17819 6307
rect 20453 6273 20487 6307
rect 22109 6273 22143 6307
rect 22661 6273 22695 6307
rect 23940 6273 23974 6307
rect 25513 6273 25547 6307
rect 26255 6273 26289 6307
rect 26433 6273 26467 6307
rect 26985 6273 27019 6307
rect 27169 6273 27203 6307
rect 27353 6273 27387 6307
rect 27997 6273 28031 6307
rect 28181 6273 28215 6307
rect 28273 6273 28307 6307
rect 28411 6273 28445 6307
rect 29101 6273 29135 6307
rect 29368 6273 29402 6307
rect 30941 6273 30975 6307
rect 31125 6273 31159 6307
rect 32137 6273 32171 6307
rect 33149 6273 33183 6307
rect 34161 6273 34195 6307
rect 34437 6273 34471 6307
rect 34529 6273 34563 6307
rect 35173 6273 35207 6307
rect 35541 6273 35575 6307
rect 36369 6273 36403 6307
rect 8033 6205 8067 6239
rect 9873 6205 9907 6239
rect 12725 6205 12759 6239
rect 18429 6205 18463 6239
rect 20729 6205 20763 6239
rect 23673 6205 23707 6239
rect 32505 6205 32539 6239
rect 7389 6137 7423 6171
rect 9137 6137 9171 6171
rect 25053 6137 25087 6171
rect 26249 6137 26283 6171
rect 32965 6137 32999 6171
rect 5641 6069 5675 6103
rect 8401 6069 8435 6103
rect 12265 6069 12299 6103
rect 14105 6069 14139 6103
rect 14933 6069 14967 6103
rect 16957 6069 16991 6103
rect 17601 6069 17635 6103
rect 21925 6069 21959 6103
rect 25697 6069 25731 6103
rect 27537 6069 27571 6103
rect 28549 6069 28583 6103
rect 30941 6069 30975 6103
rect 5089 5865 5123 5899
rect 13001 5865 13035 5899
rect 13461 5865 13495 5899
rect 14933 5865 14967 5899
rect 15117 5865 15151 5899
rect 17601 5865 17635 5899
rect 21925 5865 21959 5899
rect 26065 5865 26099 5899
rect 27905 5865 27939 5899
rect 36093 5865 36127 5899
rect 37197 5865 37231 5899
rect 5733 5797 5767 5831
rect 16037 5797 16071 5831
rect 16957 5797 16991 5831
rect 17049 5797 17083 5831
rect 19441 5797 19475 5831
rect 33517 5797 33551 5831
rect 36553 5797 36587 5831
rect 8309 5729 8343 5763
rect 14749 5729 14783 5763
rect 20545 5729 20579 5763
rect 22569 5729 22603 5763
rect 22845 5729 22879 5763
rect 29837 5729 29871 5763
rect 34713 5729 34747 5763
rect 5273 5661 5307 5695
rect 5917 5661 5951 5695
rect 6561 5661 6595 5695
rect 7481 5661 7515 5695
rect 8033 5661 8067 5695
rect 8125 5661 8159 5695
rect 8953 5661 8987 5695
rect 10793 5661 10827 5695
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 14657 5661 14691 5695
rect 14933 5661 14967 5695
rect 15853 5661 15887 5695
rect 16037 5661 16071 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 19257 5661 19291 5695
rect 19533 5661 19567 5695
rect 19809 5661 19843 5695
rect 20085 5661 20119 5695
rect 24685 5661 24719 5695
rect 26525 5661 26559 5695
rect 28549 5661 28583 5695
rect 31677 5661 31711 5695
rect 31861 5661 31895 5695
rect 33701 5661 33735 5695
rect 36737 5637 36771 5671
rect 37381 5661 37415 5695
rect 38025 5661 38059 5695
rect 9198 5593 9232 5627
rect 11060 5593 11094 5627
rect 16589 5593 16623 5627
rect 20812 5593 20846 5627
rect 24952 5593 24986 5627
rect 26770 5593 26804 5627
rect 30104 5593 30138 5627
rect 32689 5593 32723 5627
rect 32873 5593 32907 5627
rect 33057 5593 33091 5627
rect 34980 5593 35014 5627
rect 6377 5525 6411 5559
rect 7297 5525 7331 5559
rect 10333 5525 10367 5559
rect 12173 5525 12207 5559
rect 18613 5525 18647 5559
rect 28365 5525 28399 5559
rect 31217 5525 31251 5559
rect 31769 5525 31803 5559
rect 37841 5525 37875 5559
rect 4169 5321 4203 5355
rect 8769 5321 8803 5355
rect 12909 5321 12943 5355
rect 13369 5321 13403 5355
rect 15761 5321 15795 5355
rect 18153 5321 18187 5355
rect 25053 5321 25087 5355
rect 26433 5321 26467 5355
rect 28641 5321 28675 5355
rect 34253 5321 34287 5355
rect 36093 5321 36127 5355
rect 8493 5253 8527 5287
rect 9413 5253 9447 5287
rect 10425 5253 10459 5287
rect 10517 5253 10551 5287
rect 21925 5253 21959 5287
rect 26249 5253 26283 5287
rect 34069 5253 34103 5287
rect 34980 5253 35014 5287
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 6633 5185 6667 5219
rect 8217 5185 8251 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 9249 5185 9283 5219
rect 9501 5185 9535 5219
rect 9597 5185 9631 5219
rect 10241 5185 10275 5219
rect 10609 5185 10643 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12081 5185 12115 5219
rect 12541 5185 12575 5219
rect 12725 5185 12759 5219
rect 13553 5185 13587 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 14381 5185 14415 5219
rect 14648 5185 14682 5219
rect 16773 5185 16807 5219
rect 17040 5185 17074 5219
rect 18797 5185 18831 5219
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 20177 5185 20211 5219
rect 20361 5185 20395 5219
rect 21005 5185 21039 5219
rect 22109 5185 22143 5219
rect 22293 5185 22327 5219
rect 23305 5185 23339 5219
rect 23397 5185 23431 5219
rect 23673 5185 23707 5219
rect 24225 5185 24259 5219
rect 24869 5185 24903 5219
rect 26065 5185 26099 5219
rect 27261 5185 27295 5219
rect 27528 5185 27562 5219
rect 29285 5185 29319 5219
rect 30389 5185 30423 5219
rect 30573 5185 30607 5219
rect 30849 5185 30883 5219
rect 30941 5185 30975 5219
rect 32781 5185 32815 5219
rect 32873 5185 32907 5219
rect 33149 5185 33183 5219
rect 33885 5185 33919 5219
rect 34713 5185 34747 5219
rect 36737 5185 36771 5219
rect 37841 5185 37875 5219
rect 4721 5117 4755 5151
rect 33057 5117 33091 5151
rect 11989 5049 12023 5083
rect 13829 5049 13863 5083
rect 18797 5049 18831 5083
rect 20177 5049 20211 5083
rect 23121 5049 23155 5083
rect 24409 5049 24443 5083
rect 30665 5049 30699 5083
rect 32597 5049 32631 5083
rect 3801 4981 3835 5015
rect 4997 4981 5031 5015
rect 5641 4981 5675 5015
rect 7757 4981 7791 5015
rect 9781 4981 9815 5015
rect 10793 4981 10827 5015
rect 11529 4981 11563 5015
rect 19441 4981 19475 5015
rect 20821 4981 20855 5015
rect 23581 4981 23615 5015
rect 29101 4981 29135 5015
rect 36553 4981 36587 5015
rect 38025 4981 38059 5015
rect 8217 4777 8251 4811
rect 9781 4777 9815 4811
rect 10517 4777 10551 4811
rect 12449 4777 12483 4811
rect 12817 4777 12851 4811
rect 16221 4777 16255 4811
rect 16957 4777 16991 4811
rect 20637 4777 20671 4811
rect 23857 4777 23891 4811
rect 26709 4777 26743 4811
rect 28181 4777 28215 4811
rect 33609 4777 33643 4811
rect 35173 4777 35207 4811
rect 4261 4709 4295 4743
rect 13553 4709 13587 4743
rect 17877 4709 17911 4743
rect 26249 4709 26283 4743
rect 36277 4709 36311 4743
rect 6837 4641 6871 4675
rect 9413 4641 9447 4675
rect 17325 4641 17359 4675
rect 17417 4641 17451 4675
rect 19257 4641 19291 4675
rect 22477 4641 22511 4675
rect 24777 4641 24811 4675
rect 1593 4573 1627 4607
rect 3249 4573 3283 4607
rect 4445 4573 4479 4607
rect 5089 4573 5123 4607
rect 5733 4573 5767 4607
rect 6377 4573 6411 4607
rect 7104 4573 7138 4607
rect 9597 4573 9631 4607
rect 10425 4573 10459 4607
rect 10517 4573 10551 4607
rect 12541 4573 12575 4607
rect 12633 4573 12667 4607
rect 14473 4573 14507 4607
rect 14933 4573 14967 4607
rect 15209 4573 15243 4607
rect 16405 4573 16439 4607
rect 17141 4573 17175 4607
rect 18061 4573 18095 4607
rect 18521 4573 18555 4607
rect 18705 4573 18739 4607
rect 19524 4573 19558 4607
rect 21097 4573 21131 4607
rect 24593 4573 24627 4607
rect 25421 4573 25455 4607
rect 26893 4573 26927 4607
rect 27813 4573 27847 4607
rect 27997 4573 28031 4607
rect 28641 4573 28675 4607
rect 28825 4573 28859 4607
rect 29745 4573 29779 4607
rect 30389 4573 30423 4607
rect 31033 4573 31067 4607
rect 31493 4573 31527 4607
rect 31677 4573 31711 4607
rect 32229 4573 32263 4607
rect 32496 4573 32530 4607
rect 34989 4573 35023 4607
rect 35817 4573 35851 4607
rect 36461 4573 36495 4607
rect 37381 4573 37415 4607
rect 37841 4573 37875 4607
rect 10241 4505 10275 4539
rect 11161 4505 11195 4539
rect 11345 4505 11379 4539
rect 12357 4505 12391 4539
rect 13369 4505 13403 4539
rect 21281 4505 21315 4539
rect 22744 4505 22778 4539
rect 24409 4505 24443 4539
rect 25881 4505 25915 4539
rect 26065 4505 26099 4539
rect 34805 4505 34839 4539
rect 1409 4437 1443 4471
rect 3065 4437 3099 4471
rect 4905 4437 4939 4471
rect 5549 4437 5583 4471
rect 6193 4437 6227 4471
rect 10701 4437 10735 4471
rect 11529 4437 11563 4471
rect 14289 4437 14323 4471
rect 18613 4437 18647 4471
rect 21465 4437 21499 4471
rect 25237 4437 25271 4471
rect 28733 4437 28767 4471
rect 29561 4437 29595 4471
rect 30205 4437 30239 4471
rect 30849 4437 30883 4471
rect 31585 4437 31619 4471
rect 35633 4437 35667 4471
rect 37197 4437 37231 4471
rect 38025 4437 38059 4471
rect 3433 4233 3467 4267
rect 5641 4233 5675 4267
rect 21189 4233 21223 4267
rect 25881 4233 25915 4267
rect 28733 4233 28767 4267
rect 7113 4165 7147 4199
rect 11989 4165 12023 4199
rect 12817 4165 12851 4199
rect 22753 4165 22787 4199
rect 26985 4165 27019 4199
rect 27169 4165 27203 4199
rect 1593 4097 1627 4131
rect 2605 4097 2639 4131
rect 3065 4097 3099 4131
rect 3893 4097 3927 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 5825 4097 5859 4131
rect 6929 4097 6963 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 8953 4097 8987 4131
rect 9580 4097 9614 4131
rect 9719 4097 9753 4131
rect 9965 4097 9999 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 10977 4097 11011 4131
rect 12173 4097 12207 4131
rect 12633 4097 12667 4131
rect 12917 4097 12951 4131
rect 13047 4097 13081 4131
rect 13829 4097 13863 4131
rect 16129 4097 16163 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 16953 4097 16987 4131
rect 17049 4097 17083 4131
rect 18061 4097 18095 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 19165 4097 19199 4131
rect 19349 4097 19383 4131
rect 20177 4097 20211 4131
rect 20913 4097 20947 4131
rect 21097 4097 21131 4131
rect 22017 4097 22051 4131
rect 22201 4097 22235 4131
rect 22937 4097 22971 4131
rect 23029 4097 23063 4131
rect 23305 4097 23339 4131
rect 23949 4097 23983 4131
rect 24133 4097 24167 4131
rect 25237 4097 25271 4131
rect 26065 4097 26099 4131
rect 26157 4097 26191 4131
rect 26433 4097 26467 4131
rect 27353 4097 27387 4131
rect 27813 4097 27847 4131
rect 27997 4097 28031 4131
rect 28181 4097 28215 4131
rect 28917 4097 28951 4131
rect 29009 4097 29043 4131
rect 29285 4097 29319 4131
rect 29929 4097 29963 4131
rect 30665 4097 30699 4131
rect 30849 4097 30883 4131
rect 31217 4097 31251 4131
rect 32137 4097 32171 4131
rect 32321 4097 32355 4131
rect 32413 4097 32447 4131
rect 32689 4097 32723 4131
rect 33517 4097 33551 4131
rect 33977 4097 34011 4131
rect 34161 4097 34195 4131
rect 34989 4097 35023 4131
rect 35081 4097 35115 4131
rect 35725 4097 35759 4131
rect 36645 4097 36679 4131
rect 37841 4097 37875 4131
rect 7849 4029 7883 4063
rect 10885 4029 10919 4063
rect 13645 4029 13679 4063
rect 14657 4029 14691 4063
rect 14933 4029 14967 4063
rect 21833 4029 21867 4063
rect 23765 4029 23799 4063
rect 25053 4029 25087 4063
rect 30941 4029 30975 4063
rect 31033 4029 31067 4063
rect 32505 4029 32539 4063
rect 35265 4029 35299 4063
rect 2421 3961 2455 3995
rect 2881 3961 2915 3995
rect 9873 3961 9907 3995
rect 18521 3961 18555 3995
rect 25421 3961 25455 3995
rect 36461 3961 36495 3995
rect 1409 3893 1443 3927
rect 3709 3893 3743 3927
rect 4353 3893 4387 3927
rect 4997 3893 5031 3927
rect 7297 3893 7331 3927
rect 7757 3893 7791 3927
rect 8217 3893 8251 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 10425 3893 10459 3927
rect 13185 3893 13219 3927
rect 14013 3893 14047 3927
rect 15945 3893 15979 3927
rect 17233 3893 17267 3927
rect 17877 3893 17911 3927
rect 19165 3893 19199 3927
rect 20361 3893 20395 3927
rect 23213 3893 23247 3927
rect 26341 3893 26375 3927
rect 29193 3893 29227 3927
rect 29745 3893 29779 3927
rect 31401 3893 31435 3927
rect 32873 3893 32907 3927
rect 33333 3893 33367 3927
rect 33977 3893 34011 3927
rect 35909 3893 35943 3927
rect 38025 3893 38059 3927
rect 2237 3689 2271 3723
rect 7389 3689 7423 3723
rect 10333 3689 10367 3723
rect 12817 3689 12851 3723
rect 15853 3689 15887 3723
rect 18613 3689 18647 3723
rect 21557 3689 21591 3723
rect 23489 3689 23523 3723
rect 24777 3689 24811 3723
rect 26801 3689 26835 3723
rect 29009 3689 29043 3723
rect 29929 3689 29963 3723
rect 35909 3689 35943 3723
rect 1777 3621 1811 3655
rect 3065 3621 3099 3655
rect 4905 3621 4939 3655
rect 7849 3621 7883 3655
rect 10793 3621 10827 3655
rect 13277 3621 13311 3655
rect 34161 3621 34195 3655
rect 19257 3553 19291 3587
rect 22109 3553 22143 3587
rect 24409 3553 24443 3587
rect 29561 3553 29595 3587
rect 32965 3553 32999 3587
rect 33793 3553 33827 3587
rect 34713 3553 34747 3587
rect 35541 3553 35575 3587
rect 1961 3485 1995 3519
rect 2421 3485 2455 3519
rect 2789 3485 2823 3519
rect 3249 3485 3283 3519
rect 4445 3485 4479 3519
rect 5089 3485 5123 3519
rect 5549 3485 5583 3519
rect 7573 3485 7607 3519
rect 7665 3485 7699 3519
rect 7895 3485 7929 3519
rect 8953 3485 8987 3519
rect 9209 3485 9243 3519
rect 10977 3485 11011 3519
rect 11437 3485 11471 3519
rect 13461 3485 13495 3519
rect 14473 3485 14507 3519
rect 16405 3485 16439 3519
rect 16661 3485 16695 3519
rect 18245 3485 18279 3519
rect 18429 3485 18463 3519
rect 19513 3485 19547 3519
rect 21281 3485 21315 3519
rect 21373 3485 21407 3519
rect 22376 3485 22410 3519
rect 24593 3485 24627 3519
rect 25421 3485 25455 3519
rect 27636 3485 27670 3519
rect 29745 3485 29779 3519
rect 30757 3485 30791 3519
rect 32597 3485 32631 3519
rect 32781 3485 32815 3519
rect 32873 3485 32907 3519
rect 33149 3485 33183 3519
rect 33977 3485 34011 3519
rect 34897 3485 34931 3519
rect 35725 3485 35759 3519
rect 36369 3485 36403 3519
rect 37657 3485 37691 3519
rect 5794 3417 5828 3451
rect 11704 3417 11738 3451
rect 14740 3417 14774 3451
rect 25688 3417 25722 3451
rect 27885 3417 27919 3451
rect 31024 3417 31058 3451
rect 33333 3417 33367 3451
rect 4261 3349 4295 3383
rect 6929 3349 6963 3383
rect 17785 3349 17819 3383
rect 20637 3349 20671 3383
rect 32137 3349 32171 3383
rect 35081 3349 35115 3383
rect 36553 3349 36587 3383
rect 37841 3349 37875 3383
rect 2079 3145 2113 3179
rect 3065 3145 3099 3179
rect 4353 3145 4387 3179
rect 5641 3145 5675 3179
rect 10977 3145 11011 3179
rect 14197 3145 14231 3179
rect 18061 3145 18095 3179
rect 19993 3145 20027 3179
rect 21281 3145 21315 3179
rect 22063 3145 22097 3179
rect 23489 3145 23523 3179
rect 26341 3145 26375 3179
rect 1869 3077 1903 3111
rect 6644 3077 6678 3111
rect 13921 3077 13955 3111
rect 14933 3077 14967 3111
rect 16948 3077 16982 3111
rect 28457 3077 28491 3111
rect 29285 3077 29319 3111
rect 3249 3009 3283 3043
rect 3893 3009 3927 3043
rect 4537 3009 4571 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 8401 3009 8435 3043
rect 8553 3009 8587 3043
rect 8769 3009 8803 3043
rect 9597 3009 9631 3043
rect 9864 3009 9898 3043
rect 11805 3009 11839 3043
rect 12072 3009 12106 3043
rect 13645 3009 13679 3043
rect 13829 3009 13863 3043
rect 14013 3009 14047 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 15025 3009 15059 3043
rect 15761 3009 15795 3043
rect 15853 3009 15887 3043
rect 16681 3009 16715 3043
rect 18521 3009 18555 3043
rect 19717 3009 19751 3043
rect 21005 3009 21039 3043
rect 21097 3009 21131 3043
rect 23213 3009 23247 3043
rect 23305 3009 23339 3043
rect 24133 3009 24167 3043
rect 24869 3009 24903 3043
rect 25145 3009 25179 3043
rect 26249 3009 26283 3043
rect 27445 3009 27479 3043
rect 28273 3009 28307 3043
rect 29101 3009 29135 3043
rect 29745 3009 29779 3043
rect 30849 3009 30883 3043
rect 31033 3009 31067 3043
rect 31125 3009 31159 3043
rect 31401 3009 31435 3043
rect 32413 3009 32447 3043
rect 32680 3009 32714 3043
rect 34437 3009 34471 3043
rect 34989 3009 35023 3043
rect 35081 3009 35115 3043
rect 35265 3009 35299 3043
rect 35909 3009 35943 3043
rect 36093 3009 36127 3043
rect 36737 3009 36771 3043
rect 37289 3009 37323 3043
rect 19993 2941 20027 2975
rect 21833 2941 21867 2975
rect 27261 2941 27295 2975
rect 27629 2941 27663 2975
rect 28089 2941 28123 2975
rect 28917 2941 28951 2975
rect 31217 2941 31251 2975
rect 35725 2941 35759 2975
rect 2237 2873 2271 2907
rect 4997 2873 5031 2907
rect 7757 2873 7791 2907
rect 8677 2873 8711 2907
rect 15209 2873 15243 2907
rect 19809 2873 19843 2907
rect 29929 2873 29963 2907
rect 34253 2873 34287 2907
rect 2053 2805 2087 2839
rect 3709 2805 3743 2839
rect 8217 2805 8251 2839
rect 13185 2805 13219 2839
rect 16037 2805 16071 2839
rect 18705 2805 18739 2839
rect 24317 2805 24351 2839
rect 31585 2805 31619 2839
rect 33793 2805 33827 2839
rect 36553 2805 36587 2839
rect 37473 2805 37507 2839
rect 6377 2601 6411 2635
rect 8125 2601 8159 2635
rect 9321 2601 9355 2635
rect 10425 2601 10459 2635
rect 12081 2601 12115 2635
rect 14105 2601 14139 2635
rect 15853 2601 15887 2635
rect 17049 2601 17083 2635
rect 22385 2601 22419 2635
rect 26065 2601 26099 2635
rect 28825 2601 28859 2635
rect 29745 2601 29779 2635
rect 30481 2601 30515 2635
rect 32321 2601 32355 2635
rect 34897 2601 34931 2635
rect 36369 2601 36403 2635
rect 37473 2601 37507 2635
rect 2053 2533 2087 2567
rect 15393 2533 15427 2567
rect 18429 2533 18463 2567
rect 23121 2533 23155 2567
rect 27169 2533 27203 2567
rect 31217 2533 31251 2567
rect 33793 2533 33827 2567
rect 2697 2397 2731 2431
rect 3801 2397 3835 2431
rect 4721 2397 4755 2431
rect 5365 2397 5399 2431
rect 6561 2397 6595 2431
rect 7389 2397 7423 2431
rect 8309 2397 8343 2431
rect 8953 2397 8987 2431
rect 10057 2397 10091 2431
rect 12265 2397 12299 2431
rect 12725 2397 12759 2431
rect 12909 2397 12943 2431
rect 13093 2397 13127 2431
rect 14289 2397 14323 2431
rect 14841 2397 14875 2431
rect 15025 2397 15059 2431
rect 15209 2397 15243 2431
rect 16037 2397 16071 2431
rect 16681 2397 16715 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 18245 2397 18279 2431
rect 19257 2397 19291 2431
rect 19993 2397 20027 2431
rect 20729 2397 20763 2431
rect 22937 2397 22971 2431
rect 24409 2397 24443 2431
rect 25697 2397 25731 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 27721 2397 27755 2431
rect 29561 2397 29595 2431
rect 30297 2397 30331 2431
rect 31033 2397 31067 2431
rect 32137 2397 32171 2431
rect 32873 2397 32907 2431
rect 33609 2397 33643 2431
rect 34713 2397 34747 2431
rect 35449 2397 35483 2431
rect 36185 2397 36219 2431
rect 37289 2397 37323 2431
rect 1869 2329 1903 2363
rect 7021 2329 7055 2363
rect 7205 2329 7239 2363
rect 9137 2329 9171 2363
rect 10241 2329 10275 2363
rect 15117 2329 15151 2363
rect 22293 2329 22327 2363
rect 28733 2329 28767 2363
rect 2513 2261 2547 2295
rect 3985 2261 4019 2295
rect 5181 2261 5215 2295
rect 17693 2261 17727 2295
rect 19441 2261 19475 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
rect 24593 2261 24627 2295
rect 27905 2261 27939 2295
rect 33057 2261 33091 2295
rect 35633 2261 35667 2295
<< metal1 >>
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 23566 16600 23572 16652
rect 23624 16640 23630 16652
rect 23661 16643 23719 16649
rect 23661 16640 23673 16643
rect 23624 16612 23673 16640
rect 23624 16600 23630 16612
rect 23661 16609 23673 16612
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 22925 16575 22983 16581
rect 22925 16541 22937 16575
rect 22971 16572 22983 16575
rect 23014 16572 23020 16584
rect 22971 16544 23020 16572
rect 22971 16541 22983 16544
rect 22925 16535 22983 16541
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16572 23535 16575
rect 23750 16572 23756 16584
rect 23523 16544 23756 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 23400 16504 23428 16535
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 25130 16572 25136 16584
rect 25091 16544 25136 16572
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 27798 16572 27804 16584
rect 27571 16544 27804 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16572 28595 16575
rect 28810 16572 28816 16584
rect 28583 16544 28816 16572
rect 28583 16541 28595 16544
rect 28537 16535 28595 16541
rect 28810 16532 28816 16544
rect 28868 16532 28874 16584
rect 23566 16504 23572 16516
rect 23400 16476 23572 16504
rect 23566 16464 23572 16476
rect 23624 16464 23630 16516
rect 25400 16507 25458 16513
rect 25400 16473 25412 16507
rect 25446 16504 25458 16507
rect 26970 16504 26976 16516
rect 25446 16476 26976 16504
rect 25446 16473 25458 16476
rect 25400 16467 25458 16473
rect 26970 16464 26976 16476
rect 27028 16464 27034 16516
rect 28261 16507 28319 16513
rect 28261 16473 28273 16507
rect 28307 16504 28319 16507
rect 28902 16504 28908 16516
rect 28307 16476 28908 16504
rect 28307 16473 28319 16476
rect 28261 16467 28319 16473
rect 28902 16464 28908 16476
rect 28960 16464 28966 16516
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 22704 16408 22753 16436
rect 22704 16396 22710 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 23658 16436 23664 16448
rect 23619 16408 23664 16436
rect 22741 16399 22799 16405
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 26513 16439 26571 16445
rect 26513 16436 26525 16439
rect 26292 16408 26525 16436
rect 26292 16396 26298 16408
rect 26513 16405 26525 16408
rect 26559 16405 26571 16439
rect 26513 16399 26571 16405
rect 27154 16396 27160 16448
rect 27212 16436 27218 16448
rect 27341 16439 27399 16445
rect 27341 16436 27353 16439
rect 27212 16408 27353 16436
rect 27212 16396 27218 16408
rect 27341 16405 27353 16408
rect 27387 16405 27399 16439
rect 28350 16436 28356 16448
rect 28408 16445 28414 16448
rect 28317 16408 28356 16436
rect 27341 16399 27399 16405
rect 28350 16396 28356 16408
rect 28408 16399 28417 16445
rect 28445 16439 28503 16445
rect 28445 16405 28457 16439
rect 28491 16436 28503 16439
rect 29086 16436 29092 16448
rect 28491 16408 29092 16436
rect 28491 16405 28503 16408
rect 28445 16399 28503 16405
rect 28408 16396 28414 16399
rect 29086 16396 29092 16408
rect 29144 16396 29150 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 23566 16192 23572 16244
rect 23624 16232 23630 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 23624 16204 25605 16232
rect 23624 16192 23630 16204
rect 25593 16201 25605 16204
rect 25639 16201 25651 16235
rect 25593 16195 25651 16201
rect 25130 16164 25136 16176
rect 22388 16136 25136 16164
rect 22388 16105 22416 16136
rect 22646 16105 22652 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22066 16068 22385 16096
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 22066 16028 22094 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22640 16096 22652 16105
rect 22607 16068 22652 16096
rect 22373 16059 22431 16065
rect 22640 16059 22652 16068
rect 22646 16056 22652 16059
rect 22704 16056 22710 16108
rect 24228 16105 24256 16136
rect 25130 16124 25136 16136
rect 25188 16124 25194 16176
rect 26329 16167 26387 16173
rect 26329 16133 26341 16167
rect 26375 16164 26387 16167
rect 26973 16167 27031 16173
rect 26973 16164 26985 16167
rect 26375 16136 26985 16164
rect 26375 16133 26387 16136
rect 26329 16127 26387 16133
rect 26973 16133 26985 16136
rect 27019 16133 27031 16167
rect 26973 16127 27031 16133
rect 28276 16136 30236 16164
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16065 24271 16099
rect 24213 16059 24271 16065
rect 24302 16056 24308 16108
rect 24360 16096 24366 16108
rect 24469 16099 24527 16105
rect 24469 16096 24481 16099
rect 24360 16068 24481 16096
rect 24360 16056 24366 16068
rect 24469 16065 24481 16068
rect 24515 16065 24527 16099
rect 24469 16059 24527 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26234 16096 26240 16108
rect 26099 16068 26240 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26234 16056 26240 16068
rect 26292 16096 26298 16108
rect 28276 16105 28304 16136
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26292 16068 27169 16096
rect 26292 16056 26298 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27249 16099 27307 16105
rect 27249 16065 27261 16099
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 28261 16099 28319 16105
rect 28261 16065 28273 16099
rect 28307 16065 28319 16099
rect 28261 16059 28319 16065
rect 26329 16031 26387 16037
rect 26329 16028 26341 16031
rect 20772 16000 22094 16028
rect 26068 16000 26341 16028
rect 20772 15988 20778 16000
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 23532 15932 24256 15960
rect 23532 15920 23538 15932
rect 23753 15895 23811 15901
rect 23753 15861 23765 15895
rect 23799 15892 23811 15895
rect 23842 15892 23848 15904
rect 23799 15864 23848 15892
rect 23799 15861 23811 15864
rect 23753 15855 23811 15861
rect 23842 15852 23848 15864
rect 23900 15852 23906 15904
rect 24228 15892 24256 15932
rect 26068 15892 26096 16000
rect 26329 15997 26341 16000
rect 26375 15997 26387 16031
rect 26694 16028 26700 16040
rect 26329 15991 26387 15997
rect 26436 16000 26700 16028
rect 26145 15963 26203 15969
rect 26145 15929 26157 15963
rect 26191 15960 26203 15963
rect 26436 15960 26464 16000
rect 26694 15988 26700 16000
rect 26752 16028 26758 16040
rect 27264 16028 27292 16059
rect 28350 16056 28356 16108
rect 28408 16096 28414 16108
rect 28517 16099 28575 16105
rect 28517 16096 28529 16099
rect 28408 16068 28529 16096
rect 28408 16056 28414 16068
rect 28517 16065 28529 16068
rect 28563 16065 28575 16099
rect 28517 16059 28575 16065
rect 30208 16037 30236 16136
rect 30282 16056 30288 16108
rect 30340 16096 30346 16108
rect 30449 16099 30507 16105
rect 30449 16096 30461 16099
rect 30340 16068 30461 16096
rect 30340 16056 30346 16068
rect 30449 16065 30461 16068
rect 30495 16065 30507 16099
rect 30449 16059 30507 16065
rect 30742 16056 30748 16108
rect 30800 16096 30806 16108
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 30800 16068 32137 16096
rect 30800 16056 30806 16068
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 32309 16099 32367 16105
rect 32309 16065 32321 16099
rect 32355 16096 32367 16099
rect 32490 16096 32496 16108
rect 32355 16068 32496 16096
rect 32355 16065 32367 16068
rect 32309 16059 32367 16065
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 26752 16000 27292 16028
rect 30193 16031 30251 16037
rect 26752 15988 26758 16000
rect 30193 15997 30205 16031
rect 30239 15997 30251 16031
rect 30193 15991 30251 15997
rect 26970 15960 26976 15972
rect 26191 15932 26464 15960
rect 26931 15932 26976 15960
rect 26191 15929 26203 15932
rect 26145 15923 26203 15929
rect 26970 15920 26976 15932
rect 27028 15920 27034 15972
rect 28994 15892 29000 15904
rect 24228 15864 29000 15892
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 29178 15852 29184 15904
rect 29236 15892 29242 15904
rect 29641 15895 29699 15901
rect 29641 15892 29653 15895
rect 29236 15864 29653 15892
rect 29236 15852 29242 15864
rect 29641 15861 29653 15864
rect 29687 15861 29699 15895
rect 30208 15892 30236 15991
rect 31294 15892 31300 15904
rect 30208 15864 31300 15892
rect 29641 15855 29699 15861
rect 31294 15852 31300 15864
rect 31352 15852 31358 15904
rect 31570 15892 31576 15904
rect 31531 15864 31576 15892
rect 31570 15852 31576 15864
rect 31628 15852 31634 15904
rect 32122 15892 32128 15904
rect 32083 15864 32128 15892
rect 32122 15852 32128 15864
rect 32180 15852 32186 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 22833 15691 22891 15697
rect 22833 15688 22845 15691
rect 22704 15660 22845 15688
rect 22704 15648 22710 15660
rect 22833 15657 22845 15660
rect 22879 15657 22891 15691
rect 23014 15688 23020 15700
rect 22975 15660 23020 15688
rect 22833 15651 22891 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 23477 15691 23535 15697
rect 23477 15657 23489 15691
rect 23523 15688 23535 15691
rect 24302 15688 24308 15700
rect 23523 15660 24308 15688
rect 23523 15657 23535 15660
rect 23477 15651 23535 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 28902 15688 28908 15700
rect 28863 15660 28908 15688
rect 28902 15648 28908 15660
rect 28960 15648 28966 15700
rect 29917 15691 29975 15697
rect 29917 15657 29929 15691
rect 29963 15688 29975 15691
rect 30282 15688 30288 15700
rect 29963 15660 30288 15688
rect 29963 15657 29975 15660
rect 29917 15651 29975 15657
rect 30282 15648 30288 15660
rect 30340 15648 30346 15700
rect 30742 15688 30748 15700
rect 30703 15660 30748 15688
rect 30742 15648 30748 15660
rect 30800 15648 30806 15700
rect 31938 15688 31944 15700
rect 30852 15660 31944 15688
rect 28810 15620 28816 15632
rect 28771 15592 28816 15620
rect 28810 15580 28816 15592
rect 28868 15580 28874 15632
rect 30852 15620 30880 15660
rect 31938 15648 31944 15660
rect 31996 15648 32002 15700
rect 29012 15592 30880 15620
rect 29012 15564 29040 15592
rect 28994 15552 29000 15564
rect 28955 15524 29000 15552
rect 28994 15512 29000 15524
rect 29052 15512 29058 15564
rect 30837 15555 30895 15561
rect 30116 15524 30696 15552
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15484 20683 15487
rect 20714 15484 20720 15496
rect 20671 15456 20720 15484
rect 20671 15453 20683 15456
rect 20625 15447 20683 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23658 15484 23664 15496
rect 23523 15456 23664 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 20892 15419 20950 15425
rect 20892 15385 20904 15419
rect 20938 15416 20950 15419
rect 21818 15416 21824 15428
rect 20938 15388 21824 15416
rect 20938 15385 20950 15388
rect 20892 15379 20950 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 22480 15416 22508 15447
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 24581 15487 24639 15493
rect 23808 15456 23853 15484
rect 23808 15444 23814 15456
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24946 15484 24952 15496
rect 24627 15456 24952 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 25041 15487 25099 15493
rect 25041 15453 25053 15487
rect 25087 15484 25099 15487
rect 25130 15484 25136 15496
rect 25087 15456 25136 15484
rect 25087 15453 25099 15456
rect 25041 15447 25099 15453
rect 25130 15444 25136 15456
rect 25188 15484 25194 15496
rect 27154 15493 27160 15496
rect 26881 15487 26939 15493
rect 26881 15484 26893 15487
rect 25188 15456 26893 15484
rect 25188 15444 25194 15456
rect 26881 15453 26893 15456
rect 26927 15453 26939 15487
rect 27148 15484 27160 15493
rect 27115 15456 27160 15484
rect 26881 15447 26939 15453
rect 27148 15447 27160 15456
rect 27154 15444 27160 15447
rect 27212 15444 27218 15496
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15484 28779 15487
rect 29086 15484 29092 15496
rect 28767 15456 29092 15484
rect 28767 15453 28779 15456
rect 28721 15447 28779 15453
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 30116 15493 30144 15524
rect 30668 15496 30696 15524
rect 30837 15521 30849 15555
rect 30883 15552 30895 15555
rect 31110 15552 31116 15564
rect 30883 15524 31116 15552
rect 30883 15521 30895 15524
rect 30837 15515 30895 15521
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 30101 15487 30159 15493
rect 30101 15453 30113 15487
rect 30147 15453 30159 15487
rect 30101 15447 30159 15453
rect 30561 15487 30619 15493
rect 30561 15453 30573 15487
rect 30607 15453 30619 15487
rect 30561 15447 30619 15453
rect 23382 15416 23388 15428
rect 22480 15388 23388 15416
rect 23382 15376 23388 15388
rect 23440 15416 23446 15428
rect 23768 15416 23796 15444
rect 25286 15419 25344 15425
rect 25286 15416 25298 15419
rect 23440 15388 23796 15416
rect 24412 15388 25298 15416
rect 23440 15376 23446 15388
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21968 15320 22017 15348
rect 21968 15308 21974 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22830 15348 22836 15360
rect 22791 15320 22836 15348
rect 22005 15311 22063 15317
rect 22830 15308 22836 15320
rect 22888 15308 22894 15360
rect 23658 15348 23664 15360
rect 23619 15320 23664 15348
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 24412 15357 24440 15388
rect 25286 15385 25298 15388
rect 25332 15385 25344 15419
rect 29932 15416 29960 15447
rect 30466 15416 30472 15428
rect 29932 15388 30472 15416
rect 25286 15379 25344 15385
rect 30466 15376 30472 15388
rect 30524 15376 30530 15428
rect 30576 15416 30604 15447
rect 30650 15444 30656 15496
rect 30708 15484 30714 15496
rect 31294 15484 31300 15496
rect 30708 15456 30753 15484
rect 31255 15456 31300 15484
rect 30708 15444 30714 15456
rect 31294 15444 31300 15456
rect 31352 15444 31358 15496
rect 31564 15487 31622 15493
rect 31564 15453 31576 15487
rect 31610 15484 31622 15487
rect 32122 15484 32128 15496
rect 31610 15456 32128 15484
rect 31610 15453 31622 15456
rect 31564 15447 31622 15453
rect 32122 15444 32128 15456
rect 32180 15444 32186 15496
rect 30576 15388 32352 15416
rect 32324 15360 32352 15388
rect 24397 15351 24455 15357
rect 24397 15317 24409 15351
rect 24443 15317 24455 15351
rect 24397 15311 24455 15317
rect 25590 15308 25596 15360
rect 25648 15348 25654 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 25648 15320 26433 15348
rect 25648 15308 25654 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 26421 15311 26479 15317
rect 27890 15308 27896 15360
rect 27948 15348 27954 15360
rect 28261 15351 28319 15357
rect 28261 15348 28273 15351
rect 27948 15320 28273 15348
rect 27948 15308 27954 15320
rect 28261 15317 28273 15320
rect 28307 15317 28319 15351
rect 28261 15311 28319 15317
rect 32306 15308 32312 15360
rect 32364 15348 32370 15360
rect 32677 15351 32735 15357
rect 32677 15348 32689 15351
rect 32364 15320 32689 15348
rect 32364 15308 32370 15320
rect 32677 15317 32689 15320
rect 32723 15317 32735 15351
rect 32677 15311 32735 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 21818 15144 21824 15156
rect 21779 15116 21824 15144
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22741 15147 22799 15153
rect 22741 15113 22753 15147
rect 22787 15144 22799 15147
rect 22830 15144 22836 15156
rect 22787 15116 22836 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 22940 15116 23888 15144
rect 19880 15011 19938 15017
rect 19880 14977 19892 15011
rect 19926 15008 19938 15011
rect 20438 15008 20444 15020
rect 19926 14980 20444 15008
rect 19926 14977 19938 14980
rect 19880 14971 19938 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22940 15017 22968 15116
rect 23014 15036 23020 15088
rect 23072 15076 23078 15088
rect 23072 15048 23244 15076
rect 23072 15036 23078 15048
rect 23216 15017 23244 15048
rect 23860 15020 23888 15116
rect 24946 15104 24952 15156
rect 25004 15144 25010 15156
rect 25593 15147 25651 15153
rect 25593 15144 25605 15147
rect 25004 15116 25605 15144
rect 25004 15104 25010 15116
rect 25593 15113 25605 15116
rect 25639 15113 25651 15147
rect 27798 15144 27804 15156
rect 27759 15116 27804 15144
rect 25593 15107 25651 15113
rect 27798 15104 27804 15116
rect 27856 15104 27862 15156
rect 30650 15104 30656 15156
rect 30708 15144 30714 15156
rect 31389 15147 31447 15153
rect 31389 15144 31401 15147
rect 30708 15116 31401 15144
rect 30708 15104 30714 15116
rect 31389 15113 31401 15116
rect 31435 15113 31447 15147
rect 31389 15107 31447 15113
rect 25406 15076 25412 15088
rect 25367 15048 25412 15076
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 27338 15036 27344 15088
rect 27396 15076 27402 15088
rect 27617 15079 27675 15085
rect 27617 15076 27629 15079
rect 27396 15048 27629 15076
rect 27396 15036 27402 15048
rect 27617 15045 27629 15048
rect 27663 15045 27675 15079
rect 31570 15076 31576 15088
rect 27617 15039 27675 15045
rect 31128 15048 31576 15076
rect 22925 15011 22983 15017
rect 22925 14977 22937 15011
rect 22971 14977 22983 15011
rect 22925 14971 22983 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23201 14971 23259 14977
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 19628 14804 19656 14903
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 21968 14912 22293 14940
rect 21968 14900 21974 14912
rect 22281 14909 22293 14912
rect 22327 14940 22339 14943
rect 23124 14940 23152 14971
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 15008 26295 15011
rect 26418 15008 26424 15020
rect 26283 14980 26424 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 27890 14968 27896 15020
rect 27948 15008 27954 15020
rect 31128 15017 31156 15048
rect 31570 15036 31576 15048
rect 31628 15076 31634 15088
rect 32125 15079 32183 15085
rect 32125 15076 32137 15079
rect 31628 15048 32137 15076
rect 31628 15036 31634 15048
rect 32125 15045 32137 15048
rect 32171 15045 32183 15079
rect 32325 15079 32383 15085
rect 32325 15076 32337 15079
rect 32125 15039 32183 15045
rect 32232 15048 32337 15076
rect 28445 15011 28503 15017
rect 28445 15008 28457 15011
rect 27948 14980 28457 15008
rect 27948 14968 27954 14980
rect 28445 14977 28457 14980
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 31113 15011 31171 15017
rect 31113 14977 31125 15011
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 15008 31263 15011
rect 31386 15008 31392 15020
rect 31251 14980 31392 15008
rect 31251 14977 31263 14980
rect 31205 14971 31263 14977
rect 31386 14968 31392 14980
rect 31444 15008 31450 15020
rect 32232 15008 32260 15048
rect 32325 15045 32337 15048
rect 32371 15045 32383 15079
rect 32325 15039 32383 15045
rect 31444 14980 32260 15008
rect 31444 14968 31450 14980
rect 23661 14943 23719 14949
rect 23661 14940 23673 14943
rect 22327 14912 23673 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 23661 14909 23673 14912
rect 23707 14909 23719 14943
rect 23661 14903 23719 14909
rect 25041 14943 25099 14949
rect 25041 14909 25053 14943
rect 25087 14940 25099 14943
rect 26694 14940 26700 14952
rect 25087 14912 26700 14940
rect 25087 14909 25099 14912
rect 25041 14903 25099 14909
rect 26694 14900 26700 14912
rect 26752 14900 26758 14952
rect 27798 14900 27804 14952
rect 27856 14940 27862 14952
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 27856 14912 28273 14940
rect 27856 14900 27862 14912
rect 28261 14909 28273 14912
rect 28307 14909 28319 14943
rect 28261 14903 28319 14909
rect 28810 14900 28816 14952
rect 28868 14900 28874 14952
rect 26142 14872 26148 14884
rect 25424 14844 26148 14872
rect 20714 14804 20720 14816
rect 19628 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20993 14807 21051 14813
rect 20993 14773 21005 14807
rect 21039 14804 21051 14807
rect 21358 14804 21364 14816
rect 21039 14776 21364 14804
rect 21039 14773 21051 14776
rect 20993 14767 21051 14773
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 22186 14804 22192 14816
rect 22147 14776 22192 14804
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 24029 14807 24087 14813
rect 24029 14773 24041 14807
rect 24075 14804 24087 14807
rect 24394 14804 24400 14816
rect 24075 14776 24400 14804
rect 24075 14773 24087 14776
rect 24029 14767 24087 14773
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24762 14764 24768 14816
rect 24820 14804 24826 14816
rect 25424 14813 25452 14844
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 27249 14875 27307 14881
rect 27249 14841 27261 14875
rect 27295 14872 27307 14875
rect 28828 14872 28856 14900
rect 27295 14844 28856 14872
rect 27295 14841 27307 14844
rect 27249 14835 27307 14841
rect 25409 14807 25467 14813
rect 25409 14804 25421 14807
rect 24820 14776 25421 14804
rect 24820 14764 24826 14776
rect 25409 14773 25421 14776
rect 25455 14773 25467 14807
rect 26050 14804 26056 14816
rect 26011 14776 26056 14804
rect 25409 14767 25467 14773
rect 26050 14764 26056 14776
rect 26108 14764 26114 14816
rect 26160 14804 26188 14832
rect 27617 14807 27675 14813
rect 27617 14804 27629 14807
rect 26160 14776 27629 14804
rect 27617 14773 27629 14776
rect 27663 14773 27675 14807
rect 28626 14804 28632 14816
rect 28587 14776 28632 14804
rect 27617 14767 27675 14773
rect 28626 14764 28632 14776
rect 28684 14764 28690 14816
rect 32306 14804 32312 14816
rect 32267 14776 32312 14804
rect 32306 14764 32312 14776
rect 32364 14764 32370 14816
rect 32490 14804 32496 14816
rect 32451 14776 32496 14804
rect 32490 14764 32496 14776
rect 32548 14764 32554 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 18340 14572 20208 14600
rect 17586 14288 17592 14340
rect 17644 14328 17650 14340
rect 18340 14328 18368 14572
rect 18417 14535 18475 14541
rect 18417 14501 18429 14535
rect 18463 14501 18475 14535
rect 18417 14495 18475 14501
rect 18432 14464 18460 14495
rect 19705 14467 19763 14473
rect 18432 14436 19472 14464
rect 19444 14405 19472 14436
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 20070 14464 20076 14476
rect 19751 14436 20076 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20180 14464 20208 14572
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 20496 14572 20545 14600
rect 20496 14560 20502 14572
rect 20533 14569 20545 14572
rect 20579 14569 20591 14603
rect 20533 14563 20591 14569
rect 21913 14603 21971 14609
rect 21913 14569 21925 14603
rect 21959 14600 21971 14603
rect 22002 14600 22008 14612
rect 21959 14572 22008 14600
rect 21959 14569 21971 14572
rect 21913 14563 21971 14569
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 23382 14600 23388 14612
rect 23343 14572 23388 14600
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 24762 14600 24768 14612
rect 24675 14572 24768 14600
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 25406 14600 25412 14612
rect 25367 14572 25412 14600
rect 25406 14560 25412 14572
rect 25464 14560 25470 14612
rect 26694 14600 26700 14612
rect 26655 14572 26700 14600
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 27338 14600 27344 14612
rect 27299 14572 27344 14600
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 28629 14603 28687 14609
rect 28629 14569 28641 14603
rect 28675 14600 28687 14603
rect 28718 14600 28724 14612
rect 28675 14572 28724 14600
rect 28675 14569 28687 14572
rect 28629 14563 28687 14569
rect 28718 14560 28724 14572
rect 28776 14560 28782 14612
rect 30466 14560 30472 14612
rect 30524 14600 30530 14612
rect 31113 14603 31171 14609
rect 31113 14600 31125 14603
rect 30524 14572 31125 14600
rect 30524 14560 30530 14572
rect 31113 14569 31125 14572
rect 31159 14569 31171 14603
rect 31113 14563 31171 14569
rect 23290 14492 23296 14544
rect 23348 14532 23354 14544
rect 24780 14532 24808 14560
rect 25866 14532 25872 14544
rect 23348 14504 24808 14532
rect 25056 14504 25872 14532
rect 23348 14492 23354 14504
rect 20180 14436 21956 14464
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 19613 14359 19671 14365
rect 18417 14331 18475 14337
rect 18417 14328 18429 14331
rect 17644 14300 18429 14328
rect 17644 14288 17650 14300
rect 18417 14297 18429 14300
rect 18463 14297 18475 14331
rect 18708 14328 18736 14359
rect 19628 14328 19656 14359
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20548 14405 20576 14436
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 21174 14396 21180 14408
rect 21135 14368 21180 14396
rect 20533 14359 20591 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14396 21327 14399
rect 21358 14396 21364 14408
rect 21315 14368 21364 14396
rect 21315 14365 21327 14368
rect 21269 14359 21327 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 21928 14337 21956 14436
rect 25056 14408 25084 14504
rect 25866 14492 25872 14504
rect 25924 14492 25930 14544
rect 31110 14424 31116 14476
rect 31168 14464 31174 14476
rect 31205 14467 31263 14473
rect 31205 14464 31217 14467
rect 31168 14436 31217 14464
rect 31168 14424 31174 14436
rect 31205 14433 31217 14436
rect 31251 14433 31263 14467
rect 31205 14427 31263 14433
rect 22186 14396 22192 14408
rect 22099 14368 22192 14396
rect 22186 14356 22192 14368
rect 22244 14396 22250 14408
rect 23014 14396 23020 14408
rect 22244 14368 23020 14396
rect 22244 14356 22250 14368
rect 23014 14356 23020 14368
rect 23072 14356 23078 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 24302 14396 24308 14408
rect 23247 14368 24308 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 24302 14356 24308 14368
rect 24360 14356 24366 14408
rect 24397 14399 24455 14405
rect 24397 14365 24409 14399
rect 24443 14396 24455 14399
rect 25038 14396 25044 14408
rect 24443 14368 25044 14396
rect 24443 14365 24455 14368
rect 24397 14359 24455 14365
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 25590 14396 25596 14408
rect 25551 14368 25596 14396
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 25866 14396 25872 14408
rect 25827 14368 25872 14396
rect 25866 14356 25872 14368
rect 25924 14396 25930 14408
rect 26329 14399 26387 14405
rect 26329 14396 26341 14399
rect 25924 14368 26341 14396
rect 25924 14356 25930 14368
rect 26329 14365 26341 14368
rect 26375 14365 26387 14399
rect 26510 14396 26516 14408
rect 26471 14368 26516 14396
rect 26329 14359 26387 14365
rect 26510 14356 26516 14368
rect 26568 14356 26574 14408
rect 27525 14399 27583 14405
rect 27525 14365 27537 14399
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 20165 14331 20223 14337
rect 18708 14300 19748 14328
rect 18417 14291 18475 14297
rect 18598 14260 18604 14272
rect 18559 14232 18604 14260
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 19720 14260 19748 14300
rect 20165 14297 20177 14331
rect 20211 14328 20223 14331
rect 21913 14331 21971 14337
rect 20211 14300 21496 14328
rect 20211 14297 20223 14300
rect 20165 14291 20223 14297
rect 20254 14260 20260 14272
rect 19720 14232 20260 14260
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 21468 14269 21496 14300
rect 21913 14297 21925 14331
rect 21959 14297 21971 14331
rect 21913 14291 21971 14297
rect 25130 14288 25136 14340
rect 25188 14328 25194 14340
rect 25777 14331 25835 14337
rect 25777 14328 25789 14331
rect 25188 14300 25789 14328
rect 25188 14288 25194 14300
rect 25777 14297 25789 14300
rect 25823 14297 25835 14331
rect 27540 14328 27568 14359
rect 27706 14356 27712 14408
rect 27764 14396 27770 14408
rect 27801 14399 27859 14405
rect 27801 14396 27813 14399
rect 27764 14368 27813 14396
rect 27764 14356 27770 14368
rect 27801 14365 27813 14368
rect 27847 14396 27859 14399
rect 28261 14399 28319 14405
rect 28261 14396 28273 14399
rect 27847 14368 28273 14396
rect 27847 14365 27859 14368
rect 27801 14359 27859 14365
rect 28261 14365 28273 14368
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28445 14399 28503 14405
rect 28445 14365 28457 14399
rect 28491 14396 28503 14399
rect 28626 14396 28632 14408
rect 28491 14368 28632 14396
rect 28491 14365 28503 14368
rect 28445 14359 28503 14365
rect 28626 14356 28632 14368
rect 28684 14356 28690 14408
rect 29730 14396 29736 14408
rect 29691 14368 29736 14396
rect 29730 14356 29736 14368
rect 29788 14356 29794 14408
rect 30190 14396 30196 14408
rect 30151 14368 30196 14396
rect 30190 14356 30196 14368
rect 30248 14356 30254 14408
rect 30374 14396 30380 14408
rect 30335 14368 30380 14396
rect 30374 14356 30380 14368
rect 30432 14356 30438 14408
rect 30929 14399 30987 14405
rect 30929 14365 30941 14399
rect 30975 14365 30987 14399
rect 30929 14359 30987 14365
rect 31021 14399 31079 14405
rect 31021 14365 31033 14399
rect 31067 14365 31079 14399
rect 31021 14359 31079 14365
rect 27890 14328 27896 14340
rect 27540 14300 27896 14328
rect 25777 14291 25835 14297
rect 27890 14288 27896 14300
rect 27948 14288 27954 14340
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 21818 14260 21824 14272
rect 21499 14232 21824 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22097 14263 22155 14269
rect 22097 14260 22109 14263
rect 22060 14232 22109 14260
rect 22060 14220 22066 14232
rect 22097 14229 22109 14232
rect 22143 14229 22155 14263
rect 24762 14260 24768 14272
rect 24723 14232 24768 14260
rect 22097 14223 22155 14229
rect 24762 14220 24768 14232
rect 24820 14220 24826 14272
rect 24949 14263 25007 14269
rect 24949 14229 24961 14263
rect 24995 14260 25007 14263
rect 25314 14260 25320 14272
rect 24995 14232 25320 14260
rect 24995 14229 25007 14232
rect 24949 14223 25007 14229
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 27709 14263 27767 14269
rect 27709 14229 27721 14263
rect 27755 14260 27767 14263
rect 27798 14260 27804 14272
rect 27755 14232 27804 14260
rect 27755 14229 27767 14232
rect 27709 14223 27767 14229
rect 27798 14220 27804 14232
rect 27856 14220 27862 14272
rect 27982 14220 27988 14272
rect 28040 14260 28046 14272
rect 28902 14260 28908 14272
rect 28040 14232 28908 14260
rect 28040 14220 28046 14232
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 29549 14263 29607 14269
rect 29549 14260 29561 14263
rect 29052 14232 29561 14260
rect 29052 14220 29058 14232
rect 29549 14229 29561 14232
rect 29595 14229 29607 14263
rect 29549 14223 29607 14229
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 30285 14263 30343 14269
rect 30285 14260 30297 14263
rect 29696 14232 30297 14260
rect 29696 14220 29702 14232
rect 30285 14229 30297 14232
rect 30331 14229 30343 14263
rect 30944 14260 30972 14359
rect 31036 14328 31064 14359
rect 31478 14356 31484 14408
rect 31536 14396 31542 14408
rect 31665 14399 31723 14405
rect 31665 14396 31677 14399
rect 31536 14368 31677 14396
rect 31536 14356 31542 14368
rect 31665 14365 31677 14368
rect 31711 14365 31723 14399
rect 31665 14359 31723 14365
rect 31849 14399 31907 14405
rect 31849 14365 31861 14399
rect 31895 14365 31907 14399
rect 31849 14359 31907 14365
rect 31386 14328 31392 14340
rect 31036 14300 31392 14328
rect 31386 14288 31392 14300
rect 31444 14328 31450 14340
rect 31864 14328 31892 14359
rect 31444 14300 31892 14328
rect 31444 14288 31450 14300
rect 31570 14260 31576 14272
rect 30944 14232 31576 14260
rect 30285 14223 30343 14229
rect 31570 14220 31576 14232
rect 31628 14220 31634 14272
rect 31754 14260 31760 14272
rect 31715 14232 31760 14260
rect 31754 14220 31760 14232
rect 31812 14220 31818 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 18656 14028 19533 14056
rect 18656 14016 18662 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20079 14059 20137 14065
rect 20079 14025 20091 14059
rect 20125 14056 20137 14059
rect 20438 14056 20444 14068
rect 20125 14028 20444 14056
rect 20125 14025 20137 14028
rect 20079 14019 20137 14025
rect 18408 13991 18466 13997
rect 18408 13957 18420 13991
rect 18454 13988 18466 13991
rect 19242 13988 19248 14000
rect 18454 13960 19248 13988
rect 18454 13957 18466 13960
rect 18408 13951 18466 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 19536 13920 19564 14019
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 26418 14056 26424 14068
rect 26379 14028 26424 14056
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 27801 14059 27859 14065
rect 27801 14025 27813 14059
rect 27847 14056 27859 14059
rect 27982 14056 27988 14068
rect 27847 14028 27988 14056
rect 27847 14025 27859 14028
rect 27801 14019 27859 14025
rect 27982 14016 27988 14028
rect 28040 14016 28046 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 28374 14028 28549 14056
rect 28374 14000 28402 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 28902 14016 28908 14068
rect 28960 14056 28966 14068
rect 29730 14056 29736 14068
rect 28960 14028 29736 14056
rect 28960 14016 28966 14028
rect 29730 14016 29736 14028
rect 29788 14016 29794 14068
rect 31478 14056 31484 14068
rect 31439 14028 31484 14056
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 33597 14059 33655 14065
rect 33597 14025 33609 14059
rect 33643 14056 33655 14059
rect 33686 14056 33692 14068
rect 33643 14028 33692 14056
rect 33643 14025 33655 14028
rect 33597 14019 33655 14025
rect 19981 13991 20039 13997
rect 19981 13957 19993 13991
rect 20027 13988 20039 13991
rect 21358 13988 21364 14000
rect 20027 13960 21364 13988
rect 20027 13957 20039 13960
rect 19981 13951 20039 13957
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 21542 13948 21548 14000
rect 21600 13988 21606 14000
rect 21821 13991 21879 13997
rect 21821 13988 21833 13991
rect 21600 13960 21833 13988
rect 21600 13948 21606 13960
rect 21821 13957 21833 13960
rect 21867 13957 21879 13991
rect 21821 13951 21879 13957
rect 21910 13948 21916 14000
rect 21968 13988 21974 14000
rect 22021 13991 22079 13997
rect 22021 13988 22033 13991
rect 21968 13960 22033 13988
rect 21968 13948 21974 13960
rect 22021 13957 22033 13960
rect 22067 13957 22079 13991
rect 24305 13991 24363 13997
rect 24305 13988 24317 13991
rect 22021 13951 22079 13957
rect 22756 13960 24317 13988
rect 20070 13920 20076 13932
rect 19536 13892 20076 13920
rect 20070 13880 20076 13892
rect 20128 13920 20134 13932
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 20128 13892 20177 13920
rect 20128 13880 20134 13892
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17000 13824 18153 13852
rect 17000 13812 17006 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 20180 13852 20208 13883
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 21269 13923 21327 13929
rect 20312 13892 20357 13920
rect 20312 13880 20318 13892
rect 21269 13889 21281 13923
rect 21315 13920 21327 13923
rect 22370 13920 22376 13932
rect 21315 13892 22376 13920
rect 21315 13889 21327 13892
rect 21269 13883 21327 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22756 13864 22784 13960
rect 24305 13957 24317 13960
rect 24351 13957 24363 13991
rect 25590 13988 25596 14000
rect 24305 13951 24363 13957
rect 25240 13960 25596 13988
rect 24210 13920 24216 13932
rect 24171 13892 24216 13920
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24394 13920 24400 13932
rect 24355 13892 24400 13920
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 25130 13920 25136 13932
rect 25091 13892 25136 13920
rect 25130 13880 25136 13892
rect 25188 13880 25194 13932
rect 25240 13929 25268 13960
rect 25590 13948 25596 13960
rect 25648 13988 25654 14000
rect 25958 13988 25964 14000
rect 25648 13960 25964 13988
rect 25648 13948 25654 13960
rect 25958 13948 25964 13960
rect 26016 13948 26022 14000
rect 26234 13988 26240 14000
rect 26195 13960 26240 13988
rect 26234 13948 26240 13960
rect 26292 13948 26298 14000
rect 27614 13988 27620 14000
rect 27575 13960 27620 13988
rect 27614 13948 27620 13960
rect 27672 13948 27678 14000
rect 28350 13948 28356 14000
rect 28408 13948 28414 14000
rect 29086 13988 29092 14000
rect 28966 13960 29092 13988
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13920 25927 13923
rect 27706 13920 27712 13932
rect 25915 13892 27712 13920
rect 25915 13889 25927 13892
rect 25869 13883 25927 13889
rect 27706 13880 27712 13892
rect 27764 13920 27770 13932
rect 27982 13920 27988 13932
rect 27764 13892 27988 13920
rect 27764 13880 27770 13892
rect 27982 13880 27988 13892
rect 28040 13880 28046 13932
rect 28442 13920 28448 13932
rect 28403 13892 28448 13920
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 28626 13920 28632 13932
rect 28587 13892 28632 13920
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 28966 13920 28994 13960
rect 29086 13948 29092 13960
rect 29144 13948 29150 14000
rect 31294 13988 31300 14000
rect 29380 13960 31300 13988
rect 29380 13929 29408 13960
rect 31294 13948 31300 13960
rect 31352 13988 31358 14000
rect 31352 13960 31708 13988
rect 31352 13948 31358 13960
rect 31680 13932 31708 13960
rect 31754 13948 31760 14000
rect 31812 13988 31818 14000
rect 32462 13991 32520 13997
rect 32462 13988 32474 13991
rect 31812 13960 32474 13988
rect 31812 13948 31818 13960
rect 32462 13957 32474 13960
rect 32508 13957 32520 13991
rect 32462 13951 32520 13957
rect 29638 13929 29644 13932
rect 28828 13918 28994 13920
rect 28736 13892 28994 13918
rect 29365 13923 29423 13929
rect 28736 13890 28856 13892
rect 21174 13852 21180 13864
rect 20180 13824 21180 13852
rect 18141 13815 18199 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22002 13852 22008 13864
rect 21508 13824 22008 13852
rect 21508 13812 21514 13824
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 22738 13852 22744 13864
rect 22699 13824 22744 13852
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23014 13852 23020 13864
rect 22975 13824 23020 13852
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24029 13855 24087 13861
rect 24029 13852 24041 13855
rect 23716 13824 24041 13852
rect 23716 13812 23722 13824
rect 24029 13821 24041 13824
rect 24075 13852 24087 13855
rect 24486 13852 24492 13864
rect 24075 13824 24492 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 24486 13812 24492 13824
rect 24544 13812 24550 13864
rect 24581 13855 24639 13861
rect 24581 13821 24593 13855
rect 24627 13852 24639 13855
rect 24854 13852 24860 13864
rect 24627 13824 24860 13852
rect 24627 13821 24639 13824
rect 24581 13815 24639 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25409 13855 25467 13861
rect 25409 13821 25421 13855
rect 25455 13852 25467 13855
rect 26510 13852 26516 13864
rect 25455 13824 26516 13852
rect 25455 13821 25467 13824
rect 25409 13815 25467 13821
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 28261 13855 28319 13861
rect 28261 13821 28273 13855
rect 28307 13852 28319 13855
rect 28736 13852 28764 13890
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29632 13920 29644 13929
rect 29599 13892 29644 13920
rect 29365 13883 29423 13889
rect 29632 13883 29644 13892
rect 29638 13880 29644 13883
rect 29696 13880 29702 13932
rect 31202 13920 31208 13932
rect 31163 13892 31208 13920
rect 31202 13880 31208 13892
rect 31260 13920 31266 13932
rect 31260 13892 31616 13920
rect 31260 13880 31266 13892
rect 29270 13852 29276 13864
rect 28307 13824 28764 13852
rect 28966 13824 29276 13852
rect 28307 13821 28319 13824
rect 28261 13815 28319 13821
rect 19426 13744 19432 13796
rect 19484 13784 19490 13796
rect 23474 13784 23480 13796
rect 19484 13756 23480 13784
rect 19484 13744 19490 13756
rect 23474 13744 23480 13756
rect 23532 13744 23538 13796
rect 27249 13787 27307 13793
rect 27249 13753 27261 13787
rect 27295 13784 27307 13787
rect 28966 13784 28994 13824
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 30374 13812 30380 13864
rect 30432 13852 30438 13864
rect 30926 13852 30932 13864
rect 30432 13824 30932 13852
rect 30432 13812 30438 13824
rect 30926 13812 30932 13824
rect 30984 13852 30990 13864
rect 31297 13855 31355 13861
rect 31297 13852 31309 13855
rect 30984 13824 31309 13852
rect 30984 13812 30990 13824
rect 31297 13821 31309 13824
rect 31343 13821 31355 13855
rect 31481 13855 31539 13861
rect 31481 13852 31493 13855
rect 31297 13815 31355 13821
rect 31404 13824 31493 13852
rect 27295 13756 28994 13784
rect 27295 13753 27307 13756
rect 27249 13747 27307 13753
rect 31110 13744 31116 13796
rect 31168 13784 31174 13796
rect 31404 13784 31432 13824
rect 31481 13821 31493 13824
rect 31527 13821 31539 13855
rect 31588 13852 31616 13892
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32217 13923 32275 13929
rect 32217 13920 32229 13923
rect 31720 13892 32229 13920
rect 31720 13880 31726 13892
rect 32217 13889 32229 13892
rect 32263 13889 32275 13923
rect 33612 13920 33640 14019
rect 33686 14016 33692 14028
rect 33744 14016 33750 14068
rect 32217 13883 32275 13889
rect 32324 13892 33640 13920
rect 32324 13852 32352 13892
rect 31588 13824 32352 13852
rect 31481 13815 31539 13821
rect 31168 13756 31432 13784
rect 31168 13744 31174 13756
rect 21082 13716 21088 13728
rect 21043 13688 21088 13716
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 22002 13716 22008 13728
rect 21963 13688 22008 13716
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 22189 13719 22247 13725
rect 22189 13685 22201 13719
rect 22235 13716 22247 13719
rect 22278 13716 22284 13728
rect 22235 13688 22284 13716
rect 22235 13685 22247 13688
rect 22189 13679 22247 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 26142 13676 26148 13728
rect 26200 13716 26206 13728
rect 26237 13719 26295 13725
rect 26237 13716 26249 13719
rect 26200 13688 26249 13716
rect 26200 13676 26206 13688
rect 26237 13685 26249 13688
rect 26283 13716 26295 13719
rect 27617 13719 27675 13725
rect 27617 13716 27629 13719
rect 26283 13688 27629 13716
rect 26283 13685 26295 13688
rect 26237 13679 26295 13685
rect 27617 13685 27629 13688
rect 27663 13685 27675 13719
rect 27617 13679 27675 13685
rect 28813 13719 28871 13725
rect 28813 13685 28825 13719
rect 28859 13716 28871 13719
rect 29546 13716 29552 13728
rect 28859 13688 29552 13716
rect 28859 13685 28871 13688
rect 28813 13679 28871 13685
rect 29546 13676 29552 13688
rect 29604 13676 29610 13728
rect 30742 13716 30748 13728
rect 30703 13688 30748 13716
rect 30742 13676 30748 13688
rect 30800 13676 30806 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 22278 13472 22284 13524
rect 22336 13512 22342 13524
rect 23569 13515 23627 13521
rect 23569 13512 23581 13515
rect 22336 13484 23581 13512
rect 22336 13472 22342 13484
rect 23569 13481 23581 13484
rect 23615 13481 23627 13515
rect 23569 13475 23627 13481
rect 31941 13515 31999 13521
rect 31941 13481 31953 13515
rect 31987 13512 31999 13515
rect 32490 13512 32496 13524
rect 31987 13484 32496 13512
rect 31987 13481 31999 13484
rect 31941 13475 31999 13481
rect 32490 13472 32496 13484
rect 32548 13472 32554 13524
rect 20806 13444 20812 13456
rect 18524 13416 20812 13444
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 18524 13317 18552 13416
rect 20806 13404 20812 13416
rect 20864 13404 20870 13456
rect 20898 13404 20904 13456
rect 20956 13444 20962 13456
rect 21542 13444 21548 13456
rect 20956 13416 21548 13444
rect 20956 13404 20962 13416
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 29270 13404 29276 13456
rect 29328 13444 29334 13456
rect 29328 13416 29868 13444
rect 29328 13404 29334 13416
rect 29840 13388 29868 13416
rect 30742 13404 30748 13456
rect 30800 13444 30806 13456
rect 30837 13447 30895 13453
rect 30837 13444 30849 13447
rect 30800 13416 30849 13444
rect 30800 13404 30806 13416
rect 30837 13413 30849 13416
rect 30883 13413 30895 13447
rect 30837 13407 30895 13413
rect 20162 13376 20168 13388
rect 18708 13348 20168 13376
rect 18708 13317 18736 13348
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 21634 13376 21640 13388
rect 20772 13348 21640 13376
rect 20772 13336 20778 13348
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13376 23811 13379
rect 24946 13376 24952 13388
rect 23799 13348 24952 13376
rect 23799 13345 23811 13348
rect 23753 13339 23811 13345
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 26142 13376 26148 13388
rect 25056 13348 26148 13376
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 14976 13280 18061 13308
rect 14976 13268 14982 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 20070 13308 20076 13320
rect 19751 13280 20076 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 21177 13311 21235 13317
rect 21177 13277 21189 13311
rect 21223 13308 21235 13311
rect 21726 13308 21732 13320
rect 21223 13280 21732 13308
rect 21223 13277 21235 13280
rect 21177 13271 21235 13277
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 23032 13280 23489 13308
rect 19978 13200 19984 13252
rect 20036 13240 20042 13252
rect 21904 13243 21962 13249
rect 20036 13212 21128 13240
rect 20036 13200 20042 13212
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17865 13175 17923 13181
rect 17865 13172 17877 13175
rect 17184 13144 17877 13172
rect 17184 13132 17190 13144
rect 17865 13141 17877 13144
rect 17911 13141 17923 13175
rect 17865 13135 17923 13141
rect 18601 13175 18659 13181
rect 18601 13141 18613 13175
rect 18647 13172 18659 13175
rect 19334 13172 19340 13184
rect 18647 13144 19340 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 19484 13144 19809 13172
rect 19484 13132 19490 13144
rect 19797 13141 19809 13144
rect 19843 13141 19855 13175
rect 19797 13135 19855 13141
rect 20717 13175 20775 13181
rect 20717 13141 20729 13175
rect 20763 13172 20775 13175
rect 20990 13172 20996 13184
rect 20763 13144 20996 13172
rect 20763 13141 20775 13144
rect 20717 13135 20775 13141
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 21100 13181 21128 13212
rect 21904 13209 21916 13243
rect 21950 13240 21962 13243
rect 22922 13240 22928 13252
rect 21950 13212 22928 13240
rect 21950 13209 21962 13212
rect 21904 13203 21962 13209
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 21085 13175 21143 13181
rect 21085 13141 21097 13175
rect 21131 13172 21143 13175
rect 22002 13172 22008 13184
rect 21131 13144 22008 13172
rect 21131 13141 21143 13144
rect 21085 13135 21143 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 23032 13181 23060 13280
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 24854 13308 24860 13320
rect 24815 13280 24860 13308
rect 23477 13271 23535 13277
rect 24854 13268 24860 13280
rect 24912 13308 24918 13320
rect 25056 13308 25084 13348
rect 26142 13336 26148 13348
rect 26200 13376 26206 13388
rect 29546 13376 29552 13388
rect 26200 13348 26464 13376
rect 29507 13348 29552 13376
rect 26200 13336 26206 13348
rect 26436 13317 26464 13348
rect 29546 13336 29552 13348
rect 29604 13336 29610 13388
rect 29822 13376 29828 13388
rect 29735 13348 29828 13376
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 31938 13336 31944 13388
rect 31996 13376 32002 13388
rect 32125 13379 32183 13385
rect 32125 13376 32137 13379
rect 31996 13348 32137 13376
rect 31996 13336 32002 13348
rect 32125 13345 32137 13348
rect 32171 13345 32183 13379
rect 32125 13339 32183 13345
rect 24912 13280 25084 13308
rect 25133 13311 25191 13317
rect 24912 13268 24918 13280
rect 25133 13277 25145 13311
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13277 26479 13311
rect 26421 13271 26479 13277
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 25148 13240 25176 13271
rect 26510 13268 26516 13320
rect 26568 13308 26574 13320
rect 27522 13308 27528 13320
rect 26568 13280 26613 13308
rect 27483 13280 27528 13308
rect 26568 13268 26574 13280
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 27792 13311 27850 13317
rect 27792 13277 27804 13311
rect 27838 13308 27850 13311
rect 28994 13308 29000 13320
rect 27838 13280 29000 13308
rect 27838 13277 27850 13280
rect 27792 13271 27850 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 25096 13212 25176 13240
rect 26145 13243 26203 13249
rect 25096 13200 25102 13212
rect 26145 13209 26157 13243
rect 26191 13240 26203 13243
rect 29564 13240 29592 13336
rect 31021 13311 31079 13317
rect 31021 13277 31033 13311
rect 31067 13308 31079 13311
rect 31202 13308 31208 13320
rect 31067 13280 31208 13308
rect 31067 13277 31079 13280
rect 31021 13271 31079 13277
rect 31202 13268 31208 13280
rect 31260 13268 31266 13320
rect 31849 13311 31907 13317
rect 31849 13277 31861 13311
rect 31895 13308 31907 13311
rect 32398 13308 32404 13320
rect 31895 13280 32404 13308
rect 31895 13277 31907 13280
rect 31849 13271 31907 13277
rect 32398 13268 32404 13280
rect 32456 13268 32462 13320
rect 30282 13240 30288 13252
rect 26191 13212 26464 13240
rect 29564 13212 30288 13240
rect 26191 13209 26203 13212
rect 26145 13203 26203 13209
rect 26436 13184 26464 13212
rect 30282 13200 30288 13212
rect 30340 13240 30346 13252
rect 31113 13243 31171 13249
rect 31113 13240 31125 13243
rect 30340 13212 31125 13240
rect 30340 13200 30346 13212
rect 31113 13209 31125 13212
rect 31159 13209 31171 13243
rect 31113 13203 31171 13209
rect 23017 13175 23075 13181
rect 23017 13172 23029 13175
rect 22152 13144 23029 13172
rect 22152 13132 22158 13144
rect 23017 13141 23029 13144
rect 23063 13141 23075 13175
rect 23750 13172 23756 13184
rect 23711 13144 23756 13172
rect 23017 13135 23075 13141
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 26326 13172 26332 13184
rect 26287 13144 26332 13172
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 26418 13132 26424 13184
rect 26476 13132 26482 13184
rect 26697 13175 26755 13181
rect 26697 13141 26709 13175
rect 26743 13172 26755 13175
rect 27338 13172 27344 13184
rect 26743 13144 27344 13172
rect 26743 13141 26755 13144
rect 26697 13135 26755 13141
rect 27338 13132 27344 13144
rect 27396 13132 27402 13184
rect 28442 13132 28448 13184
rect 28500 13172 28506 13184
rect 28718 13172 28724 13184
rect 28500 13144 28724 13172
rect 28500 13132 28506 13144
rect 28718 13132 28724 13144
rect 28776 13172 28782 13184
rect 28905 13175 28963 13181
rect 28905 13172 28917 13175
rect 28776 13144 28917 13172
rect 28776 13132 28782 13144
rect 28905 13141 28917 13144
rect 28951 13141 28963 13175
rect 28905 13135 28963 13141
rect 31202 13132 31208 13184
rect 31260 13172 31266 13184
rect 31386 13172 31392 13184
rect 31260 13144 31305 13172
rect 31347 13144 31392 13172
rect 31260 13132 31266 13144
rect 31386 13132 31392 13144
rect 31444 13132 31450 13184
rect 31478 13132 31484 13184
rect 31536 13172 31542 13184
rect 32125 13175 32183 13181
rect 32125 13172 32137 13175
rect 31536 13144 32137 13172
rect 31536 13132 31542 13144
rect 32125 13141 32137 13144
rect 32171 13141 32183 13175
rect 32125 13135 32183 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 21048 12940 22201 12968
rect 21048 12928 21054 12940
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22370 12968 22376 12980
rect 22331 12940 22376 12968
rect 22189 12931 22247 12937
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24578 12968 24584 12980
rect 24268 12940 24584 12968
rect 24268 12928 24274 12940
rect 24578 12928 24584 12940
rect 24636 12968 24642 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24636 12940 24685 12968
rect 24636 12928 24642 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 24673 12931 24731 12937
rect 25133 12971 25191 12977
rect 25133 12937 25145 12971
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 25869 12971 25927 12977
rect 25869 12937 25881 12971
rect 25915 12968 25927 12971
rect 26234 12968 26240 12980
rect 25915 12940 26240 12968
rect 25915 12937 25927 12940
rect 25869 12931 25927 12937
rect 19242 12900 19248 12912
rect 19203 12872 19248 12900
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 23560 12903 23618 12909
rect 23560 12869 23572 12903
rect 23606 12900 23618 12903
rect 25148 12900 25176 12931
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 27614 12928 27620 12980
rect 27672 12968 27678 12980
rect 28629 12971 28687 12977
rect 28629 12968 28641 12971
rect 27672 12940 28641 12968
rect 27672 12928 27678 12940
rect 28629 12937 28641 12940
rect 28675 12937 28687 12971
rect 30926 12968 30932 12980
rect 28629 12931 28687 12937
rect 29932 12940 30788 12968
rect 30887 12940 30932 12968
rect 23606 12872 25176 12900
rect 25415 12872 29316 12900
rect 23606 12869 23618 12872
rect 23560 12863 23618 12869
rect 9674 12792 9680 12844
rect 9732 12841 9738 12844
rect 9732 12832 9743 12841
rect 10502 12832 10508 12844
rect 9732 12804 9777 12832
rect 10463 12804 10508 12832
rect 9732 12795 9743 12804
rect 9732 12792 9738 12795
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17678 12832 17684 12844
rect 17635 12804 17684 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17420 12764 17448 12795
rect 17678 12792 17684 12804
rect 17736 12832 17742 12844
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 17736 12804 18153 12832
rect 17736 12792 17742 12804
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 19426 12832 19432 12844
rect 18141 12795 18199 12801
rect 18432 12804 19432 12832
rect 18432 12773 18460 12804
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 19978 12832 19984 12844
rect 19935 12804 19984 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 21634 12792 21640 12844
rect 21692 12832 21698 12844
rect 23293 12835 23351 12841
rect 23293 12832 23305 12835
rect 21692 12804 23305 12832
rect 21692 12792 21698 12804
rect 23293 12801 23305 12804
rect 23339 12801 23351 12835
rect 25314 12832 25320 12844
rect 25275 12804 25320 12832
rect 23293 12795 23351 12801
rect 25314 12792 25320 12804
rect 25372 12792 25378 12844
rect 18417 12767 18475 12773
rect 17420 12736 17632 12764
rect 17604 12708 17632 12736
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 18923 12736 20177 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 20165 12733 20177 12736
rect 20211 12764 20223 12767
rect 20254 12764 20260 12776
rect 20211 12736 20260 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21821 12767 21879 12773
rect 21821 12733 21833 12767
rect 21867 12764 21879 12767
rect 22278 12764 22284 12776
rect 21867 12736 22284 12764
rect 21867 12733 21879 12736
rect 21821 12727 21879 12733
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 17586 12656 17592 12708
rect 17644 12656 17650 12708
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 18325 12699 18383 12705
rect 18325 12696 18337 12699
rect 18012 12668 18337 12696
rect 18012 12656 18018 12668
rect 18325 12665 18337 12668
rect 18371 12665 18383 12699
rect 18325 12659 18383 12665
rect 19260 12668 22232 12696
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 11606 12628 11612 12640
rect 10367 12600 11612 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 17402 12628 17408 12640
rect 17363 12600 17408 12628
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19260 12637 19288 12668
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 19208 12600 19257 12628
rect 19208 12588 19214 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19245 12591 19303 12597
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12628 19487 12631
rect 20806 12628 20812 12640
rect 19475 12600 20812 12628
rect 19475 12597 19487 12600
rect 19429 12591 19487 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 22204 12637 22232 12668
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22646 12628 22652 12640
rect 22235 12600 22652 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22646 12588 22652 12600
rect 22704 12628 22710 12640
rect 25415 12628 25443 12872
rect 26142 12832 26148 12844
rect 26103 12804 26148 12832
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12832 26295 12835
rect 26418 12832 26424 12844
rect 26283 12804 26424 12832
rect 26283 12801 26295 12804
rect 26237 12795 26295 12801
rect 26418 12792 26424 12804
rect 26476 12832 26482 12844
rect 26970 12832 26976 12844
rect 26476 12804 26976 12832
rect 26476 12792 26482 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27338 12832 27344 12844
rect 27251 12804 27344 12832
rect 27338 12792 27344 12804
rect 27396 12832 27402 12844
rect 27396 12804 28396 12832
rect 27396 12792 27402 12804
rect 28368 12776 28396 12804
rect 28626 12792 28632 12844
rect 28684 12832 28690 12844
rect 28813 12835 28871 12841
rect 28813 12832 28825 12835
rect 28684 12804 28825 12832
rect 28684 12792 28690 12804
rect 28813 12801 28825 12804
rect 28859 12801 28871 12835
rect 28994 12832 29000 12844
rect 28955 12804 29000 12832
rect 28813 12795 28871 12801
rect 28994 12792 29000 12804
rect 29052 12792 29058 12844
rect 26053 12767 26111 12773
rect 26053 12733 26065 12767
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 26068 12696 26096 12727
rect 26326 12724 26332 12776
rect 26384 12764 26390 12776
rect 26878 12764 26884 12776
rect 26384 12736 26884 12764
rect 26384 12724 26390 12736
rect 26878 12724 26884 12736
rect 26936 12724 26942 12776
rect 27617 12767 27675 12773
rect 27617 12733 27629 12767
rect 27663 12764 27675 12767
rect 27982 12764 27988 12776
rect 27663 12736 27988 12764
rect 27663 12733 27675 12736
rect 27617 12727 27675 12733
rect 27982 12724 27988 12736
rect 28040 12724 28046 12776
rect 28350 12724 28356 12776
rect 28408 12764 28414 12776
rect 28905 12767 28963 12773
rect 28905 12764 28917 12767
rect 28408 12736 28917 12764
rect 28408 12724 28414 12736
rect 28905 12733 28917 12736
rect 28951 12733 28963 12767
rect 28905 12727 28963 12733
rect 29089 12767 29147 12773
rect 29089 12733 29101 12767
rect 29135 12733 29147 12767
rect 29288 12764 29316 12872
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 29932 12841 29960 12940
rect 30561 12903 30619 12909
rect 30561 12869 30573 12903
rect 30607 12900 30619 12903
rect 30650 12900 30656 12912
rect 30607 12872 30656 12900
rect 30607 12869 30619 12872
rect 30561 12863 30619 12869
rect 30650 12860 30656 12872
rect 30708 12860 30714 12912
rect 30760 12909 30788 12940
rect 30926 12928 30932 12940
rect 30984 12928 30990 12980
rect 31386 12928 31392 12980
rect 31444 12968 31450 12980
rect 32493 12971 32551 12977
rect 32493 12968 32505 12971
rect 31444 12940 32505 12968
rect 31444 12928 31450 12940
rect 32493 12937 32505 12940
rect 32539 12937 32551 12971
rect 32493 12931 32551 12937
rect 30760 12903 30835 12909
rect 30760 12872 30789 12903
rect 30777 12869 30789 12872
rect 30823 12900 30835 12903
rect 31018 12900 31024 12912
rect 30823 12872 31024 12900
rect 30823 12869 30835 12872
rect 30777 12863 30835 12869
rect 31018 12860 31024 12872
rect 31076 12900 31082 12912
rect 31202 12900 31208 12912
rect 31076 12872 31208 12900
rect 31076 12860 31082 12872
rect 31202 12860 31208 12872
rect 31260 12860 31266 12912
rect 29917 12835 29975 12841
rect 29917 12801 29929 12835
rect 29963 12801 29975 12835
rect 30668 12832 30696 12860
rect 31294 12832 31300 12844
rect 30668 12804 31300 12832
rect 29917 12795 29975 12801
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 31389 12835 31447 12841
rect 31389 12801 31401 12835
rect 31435 12832 31447 12835
rect 31478 12832 31484 12844
rect 31435 12804 31484 12832
rect 31435 12801 31447 12804
rect 31389 12795 31447 12801
rect 31478 12792 31484 12804
rect 31536 12792 31542 12844
rect 31573 12835 31631 12841
rect 31573 12801 31585 12835
rect 31619 12832 31631 12835
rect 32306 12832 32312 12844
rect 31619 12804 31754 12832
rect 32267 12804 32312 12832
rect 31619 12801 31631 12804
rect 31573 12795 31631 12801
rect 31726 12764 31754 12804
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 32398 12792 32404 12844
rect 32456 12832 32462 12844
rect 32456 12804 32501 12832
rect 32456 12792 32462 12804
rect 33134 12792 33140 12844
rect 33192 12832 33198 12844
rect 33781 12835 33839 12841
rect 33781 12832 33793 12835
rect 33192 12804 33793 12832
rect 33192 12792 33198 12804
rect 33781 12801 33793 12804
rect 33827 12801 33839 12835
rect 33781 12795 33839 12801
rect 33318 12764 33324 12776
rect 29288 12736 31515 12764
rect 31726 12736 33324 12764
rect 29089 12727 29147 12733
rect 26510 12696 26516 12708
rect 26068 12668 26516 12696
rect 26510 12656 26516 12668
rect 26568 12656 26574 12708
rect 28074 12656 28080 12708
rect 28132 12696 28138 12708
rect 28718 12696 28724 12708
rect 28132 12668 28724 12696
rect 28132 12656 28138 12668
rect 28718 12656 28724 12668
rect 28776 12696 28782 12708
rect 29104 12696 29132 12727
rect 28776 12668 29132 12696
rect 28776 12656 28782 12668
rect 22704 12600 25443 12628
rect 22704 12588 22710 12600
rect 28994 12588 29000 12640
rect 29052 12628 29058 12640
rect 29638 12628 29644 12640
rect 29052 12600 29644 12628
rect 29052 12588 29058 12600
rect 29638 12588 29644 12600
rect 29696 12588 29702 12640
rect 29914 12588 29920 12640
rect 29972 12628 29978 12640
rect 30101 12631 30159 12637
rect 30101 12628 30113 12631
rect 29972 12600 30113 12628
rect 29972 12588 29978 12600
rect 30101 12597 30113 12600
rect 30147 12597 30159 12631
rect 30101 12591 30159 12597
rect 30282 12588 30288 12640
rect 30340 12628 30346 12640
rect 30745 12631 30803 12637
rect 30745 12628 30757 12631
rect 30340 12600 30757 12628
rect 30340 12588 30346 12600
rect 30745 12597 30757 12600
rect 30791 12597 30803 12631
rect 31386 12628 31392 12640
rect 31347 12600 31392 12628
rect 30745 12591 30803 12597
rect 31386 12588 31392 12600
rect 31444 12588 31450 12640
rect 31487 12628 31515 12736
rect 33318 12724 33324 12736
rect 33376 12764 33382 12776
rect 33597 12767 33655 12773
rect 33597 12764 33609 12767
rect 33376 12736 33609 12764
rect 33376 12724 33382 12736
rect 33597 12733 33609 12736
rect 33643 12733 33655 12767
rect 33597 12727 33655 12733
rect 33689 12767 33747 12773
rect 33689 12733 33701 12767
rect 33735 12733 33747 12767
rect 33870 12764 33876 12776
rect 33831 12736 33876 12764
rect 33689 12727 33747 12733
rect 31570 12656 31576 12708
rect 31628 12696 31634 12708
rect 32125 12699 32183 12705
rect 32125 12696 32137 12699
rect 31628 12668 32137 12696
rect 31628 12656 31634 12668
rect 32125 12665 32137 12668
rect 32171 12665 32183 12699
rect 32125 12659 32183 12665
rect 33502 12656 33508 12708
rect 33560 12696 33566 12708
rect 33704 12696 33732 12727
rect 33870 12724 33876 12736
rect 33928 12724 33934 12776
rect 33560 12668 33732 12696
rect 33560 12656 33566 12668
rect 32214 12628 32220 12640
rect 31487 12600 32220 12628
rect 32214 12588 32220 12600
rect 32272 12588 32278 12640
rect 32674 12628 32680 12640
rect 32635 12600 32680 12628
rect 32674 12588 32680 12600
rect 32732 12588 32738 12640
rect 33413 12631 33471 12637
rect 33413 12597 33425 12631
rect 33459 12628 33471 12631
rect 33962 12628 33968 12640
rect 33459 12600 33968 12628
rect 33459 12597 33471 12600
rect 33413 12591 33471 12597
rect 33962 12588 33968 12600
rect 34020 12588 34026 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12424 10011 12427
rect 10502 12424 10508 12436
rect 9999 12396 10508 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 16390 12424 16396 12436
rect 16303 12396 16396 12424
rect 16390 12384 16396 12396
rect 16448 12424 16454 12436
rect 19150 12424 19156 12436
rect 16448 12396 19156 12424
rect 16448 12384 16454 12396
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 19889 12427 19947 12433
rect 19889 12393 19901 12427
rect 19935 12424 19947 12427
rect 19978 12424 19984 12436
rect 19935 12396 19984 12424
rect 19935 12393 19947 12396
rect 19889 12387 19947 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 21726 12424 21732 12436
rect 20088 12396 21732 12424
rect 18325 12359 18383 12365
rect 18325 12325 18337 12359
rect 18371 12356 18383 12359
rect 18414 12356 18420 12368
rect 18371 12328 18420 12356
rect 18371 12325 18383 12328
rect 18325 12319 18383 12325
rect 18414 12316 18420 12328
rect 18472 12356 18478 12368
rect 19337 12359 19395 12365
rect 19337 12356 19349 12359
rect 18472 12328 19349 12356
rect 18472 12316 18478 12328
rect 19337 12325 19349 12328
rect 19383 12325 19395 12359
rect 19337 12319 19395 12325
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 8294 12288 8300 12300
rect 6779 12260 8300 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 8294 12248 8300 12260
rect 8352 12288 8358 12300
rect 9490 12288 9496 12300
rect 8352 12260 9496 12288
rect 8352 12248 8358 12260
rect 9490 12248 9496 12260
rect 9548 12288 9554 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9548 12260 9597 12288
rect 9548 12248 9554 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 20088 12288 20116 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 24397 12427 24455 12433
rect 24397 12393 24409 12427
rect 24443 12424 24455 12427
rect 24762 12424 24768 12436
rect 24443 12396 24768 12424
rect 24443 12393 24455 12396
rect 24397 12387 24455 12393
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 24946 12384 24952 12436
rect 25004 12424 25010 12436
rect 28721 12427 28779 12433
rect 28721 12424 28733 12427
rect 25004 12396 28733 12424
rect 25004 12384 25010 12396
rect 28721 12393 28733 12396
rect 28767 12393 28779 12427
rect 28721 12387 28779 12393
rect 30009 12427 30067 12433
rect 30009 12393 30021 12427
rect 30055 12424 30067 12427
rect 30190 12424 30196 12436
rect 30055 12396 30196 12424
rect 30055 12393 30067 12396
rect 30009 12387 30067 12393
rect 24486 12316 24492 12368
rect 24544 12356 24550 12368
rect 24544 12328 24808 12356
rect 24544 12316 24550 12328
rect 23290 12288 23296 12300
rect 18104 12260 20116 12288
rect 23251 12260 23296 12288
rect 18104 12248 18110 12260
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 24394 12248 24400 12300
rect 24452 12288 24458 12300
rect 24780 12297 24808 12328
rect 27154 12316 27160 12368
rect 27212 12356 27218 12368
rect 27433 12359 27491 12365
rect 27433 12356 27445 12359
rect 27212 12328 27445 12356
rect 27212 12316 27218 12328
rect 27433 12325 27445 12328
rect 27479 12325 27491 12359
rect 27433 12319 27491 12325
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 24452 12260 24593 12288
rect 24452 12248 24458 12260
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 24765 12291 24823 12297
rect 24765 12257 24777 12291
rect 24811 12257 24823 12291
rect 28736 12288 28764 12387
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 30101 12291 30159 12297
rect 30101 12288 30113 12291
rect 28736 12260 30113 12288
rect 24765 12251 24823 12257
rect 30101 12257 30113 12260
rect 30147 12288 30159 12291
rect 31110 12288 31116 12300
rect 30147 12260 31116 12288
rect 30147 12257 30159 12260
rect 30101 12251 30159 12257
rect 31110 12248 31116 12260
rect 31168 12248 31174 12300
rect 6914 12220 6920 12232
rect 6875 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8570 12220 8576 12232
rect 7883 12192 8576 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9125 12183 9183 12189
rect 9140 12152 9168 12183
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 11330 12220 11336 12232
rect 11291 12192 11336 12220
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13872 12192 14565 12220
rect 13872 12180 13878 12192
rect 14553 12189 14565 12192
rect 14599 12220 14611 12223
rect 16206 12220 16212 12232
rect 14599 12192 16212 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17212 12223 17270 12229
rect 17212 12189 17224 12223
rect 17258 12220 17270 12223
rect 17258 12192 17356 12220
rect 17258 12189 17270 12192
rect 17212 12183 17270 12189
rect 9950 12152 9956 12164
rect 9140 12124 9956 12152
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 10502 12152 10508 12164
rect 10463 12124 10508 12152
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 14737 12155 14795 12161
rect 14737 12121 14749 12155
rect 14783 12152 14795 12155
rect 14826 12152 14832 12164
rect 14783 12124 14832 12152
rect 14783 12121 14795 12124
rect 14737 12115 14795 12121
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 5868 12056 7113 12084
rect 5868 12044 5874 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7101 12047 7159 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9214 12084 9220 12096
rect 8987 12056 9220 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10468 12056 10609 12084
rect 10468 12044 10474 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10744 12056 11161 12084
rect 10744 12044 10750 12056
rect 11149 12053 11161 12056
rect 11195 12053 11207 12087
rect 11149 12047 11207 12053
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12434 12084 12440 12096
rect 11931 12056 12440 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 17328 12084 17356 12192
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19208 12192 19625 12220
rect 19208 12180 19214 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12220 20683 12223
rect 20714 12220 20720 12232
rect 20671 12192 20720 12220
rect 20671 12189 20683 12192
rect 20625 12183 20683 12189
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 21358 12180 21364 12232
rect 21416 12220 21422 12232
rect 21634 12220 21640 12232
rect 21416 12192 21640 12220
rect 21416 12180 21422 12192
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 21784 12192 23029 12220
rect 21784 12180 21790 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 23017 12183 23075 12189
rect 23124 12192 24685 12220
rect 17494 12112 17500 12164
rect 17552 12152 17558 12164
rect 20070 12152 20076 12164
rect 17552 12124 20076 12152
rect 17552 12112 17558 12124
rect 20070 12112 20076 12124
rect 20128 12152 20134 12164
rect 20530 12152 20536 12164
rect 20128 12124 20536 12152
rect 20128 12112 20134 12124
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20892 12155 20950 12161
rect 20892 12121 20904 12155
rect 20938 12152 20950 12155
rect 21082 12152 21088 12164
rect 20938 12124 21088 12152
rect 20938 12121 20950 12124
rect 20892 12115 20950 12121
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21232 12124 22324 12152
rect 21232 12112 21238 12124
rect 17402 12084 17408 12096
rect 17328 12056 17408 12084
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 19484 12056 19533 12084
rect 19484 12044 19490 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 21358 12084 21364 12096
rect 19751 12056 21364 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 21542 12044 21548 12096
rect 21600 12084 21606 12096
rect 21818 12084 21824 12096
rect 21600 12056 21824 12084
rect 21600 12044 21606 12056
rect 21818 12044 21824 12056
rect 21876 12084 21882 12096
rect 22005 12087 22063 12093
rect 22005 12084 22017 12087
rect 21876 12056 22017 12084
rect 21876 12044 21882 12056
rect 22005 12053 22017 12056
rect 22051 12053 22063 12087
rect 22296 12084 22324 12124
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 22738 12152 22744 12164
rect 22428 12124 22744 12152
rect 22428 12112 22434 12124
rect 22738 12112 22744 12124
rect 22796 12152 22802 12164
rect 23124 12152 23152 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24857 12223 24915 12229
rect 24857 12189 24869 12223
rect 24903 12189 24915 12223
rect 25590 12220 25596 12232
rect 25551 12192 25596 12220
rect 24857 12183 24915 12189
rect 22796 12124 23152 12152
rect 22796 12112 22802 12124
rect 24578 12112 24584 12164
rect 24636 12152 24642 12164
rect 24872 12152 24900 12183
rect 25590 12180 25596 12192
rect 25648 12180 25654 12232
rect 27706 12220 27712 12232
rect 27667 12192 27712 12220
rect 27706 12180 27712 12192
rect 27764 12220 27770 12232
rect 27982 12220 27988 12232
rect 27764 12192 27988 12220
rect 27764 12180 27770 12192
rect 27982 12180 27988 12192
rect 28040 12180 28046 12232
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 24636 12124 24900 12152
rect 25860 12155 25918 12161
rect 24636 12112 24642 12124
rect 25860 12121 25872 12155
rect 25906 12152 25918 12155
rect 26050 12152 26056 12164
rect 25906 12124 26056 12152
rect 25906 12121 25918 12124
rect 25860 12115 25918 12121
rect 26050 12112 26056 12124
rect 26108 12112 26114 12164
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 26804 12124 27445 12152
rect 25682 12084 25688 12096
rect 22296 12056 25688 12084
rect 22005 12047 22063 12053
rect 25682 12044 25688 12056
rect 25740 12084 25746 12096
rect 26804 12084 26832 12124
rect 27433 12121 27445 12124
rect 27479 12152 27491 12155
rect 28626 12152 28632 12164
rect 27479 12124 28488 12152
rect 28587 12124 28632 12152
rect 27479 12121 27491 12124
rect 27433 12115 27491 12121
rect 26970 12084 26976 12096
rect 25740 12056 26832 12084
rect 26931 12056 26976 12084
rect 25740 12044 25746 12056
rect 26970 12044 26976 12056
rect 27028 12044 27034 12096
rect 27617 12087 27675 12093
rect 27617 12053 27629 12087
rect 27663 12084 27675 12087
rect 27798 12084 27804 12096
rect 27663 12056 27804 12084
rect 27663 12053 27675 12056
rect 27617 12047 27675 12053
rect 27798 12044 27804 12056
rect 27856 12084 27862 12096
rect 28258 12084 28264 12096
rect 27856 12056 28264 12084
rect 27856 12044 27862 12056
rect 28258 12044 28264 12056
rect 28316 12044 28322 12096
rect 28460 12084 28488 12124
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 29840 12152 29868 12183
rect 29914 12180 29920 12232
rect 29972 12220 29978 12232
rect 30742 12220 30748 12232
rect 29972 12192 30017 12220
rect 30703 12192 30748 12220
rect 29972 12180 29978 12192
rect 30742 12180 30748 12192
rect 30800 12180 30806 12232
rect 31202 12220 31208 12232
rect 31163 12192 31208 12220
rect 31202 12180 31208 12192
rect 31260 12220 31266 12232
rect 31260 12192 31708 12220
rect 31260 12180 31266 12192
rect 31680 12164 31708 12192
rect 32674 12180 32680 12232
rect 32732 12220 32738 12232
rect 33045 12223 33103 12229
rect 33045 12220 33057 12223
rect 32732 12192 33057 12220
rect 32732 12180 32738 12192
rect 33045 12189 33057 12192
rect 33091 12189 33103 12223
rect 33318 12220 33324 12232
rect 33279 12192 33324 12220
rect 33045 12183 33103 12189
rect 33318 12180 33324 12192
rect 33376 12180 33382 12232
rect 30650 12152 30656 12164
rect 29840 12124 30656 12152
rect 30650 12112 30656 12124
rect 30708 12112 30714 12164
rect 31478 12161 31484 12164
rect 31472 12115 31484 12161
rect 31536 12152 31542 12164
rect 31536 12124 31572 12152
rect 31478 12112 31484 12115
rect 31536 12112 31542 12124
rect 31662 12112 31668 12164
rect 31720 12112 31726 12164
rect 29638 12084 29644 12096
rect 28460 12056 29644 12084
rect 29638 12044 29644 12056
rect 29696 12044 29702 12096
rect 30558 12084 30564 12096
rect 30519 12056 30564 12084
rect 30558 12044 30564 12056
rect 30616 12044 30622 12096
rect 32582 12084 32588 12096
rect 32543 12056 32588 12084
rect 32582 12044 32588 12056
rect 32640 12044 32646 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 21174 11880 21180 11892
rect 12584 11852 21180 11880
rect 12584 11840 12590 11852
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 22002 11840 22008 11892
rect 22060 11880 22066 11892
rect 22097 11883 22155 11889
rect 22097 11880 22109 11883
rect 22060 11852 22109 11880
rect 22060 11840 22066 11852
rect 22097 11849 22109 11852
rect 22143 11849 22155 11883
rect 22370 11880 22376 11892
rect 22331 11852 22376 11880
rect 22097 11843 22155 11849
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 22922 11880 22928 11892
rect 22883 11852 22928 11880
rect 22922 11840 22928 11852
rect 22980 11840 22986 11892
rect 28994 11840 29000 11892
rect 29052 11880 29058 11892
rect 30193 11883 30251 11889
rect 30193 11880 30205 11883
rect 29052 11852 30205 11880
rect 29052 11840 29058 11852
rect 30193 11849 30205 11852
rect 30239 11880 30251 11883
rect 31018 11880 31024 11892
rect 30239 11852 30880 11880
rect 30979 11852 31024 11880
rect 30239 11849 30251 11852
rect 30193 11843 30251 11849
rect 7006 11812 7012 11824
rect 6380 11784 7012 11812
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 6380 11753 6408 11784
rect 7006 11772 7012 11784
rect 7064 11812 7070 11824
rect 10410 11812 10416 11824
rect 7064 11784 10416 11812
rect 7064 11772 7070 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 6365 11707 6423 11713
rect 6472 11716 6633 11744
rect 6472 11676 6500 11716
rect 6621 11713 6633 11716
rect 6667 11713 6679 11747
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 6621 11707 6679 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9140 11753 9168 11784
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11762 11815 11820 11821
rect 11762 11812 11774 11815
rect 11664 11784 11774 11812
rect 11664 11772 11670 11784
rect 11762 11781 11774 11784
rect 11808 11781 11820 11815
rect 11762 11775 11820 11781
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 16025 11815 16083 11821
rect 13320 11784 14228 11812
rect 13320 11772 13326 11784
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9381 11747 9439 11753
rect 9381 11744 9393 11747
rect 9272 11716 9393 11744
rect 9272 11704 9278 11716
rect 9381 11713 9393 11716
rect 9427 11713 9439 11747
rect 9381 11707 9439 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 12342 11744 12348 11756
rect 11563 11716 12348 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 13354 11744 13360 11756
rect 13315 11716 13360 11744
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13538 11744 13544 11756
rect 13499 11716 13544 11744
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13998 11744 14004 11756
rect 13959 11716 14004 11744
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14200 11753 14228 11784
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 17190 11815 17248 11821
rect 17190 11812 17202 11815
rect 16071 11784 17202 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 17190 11781 17202 11784
rect 17236 11781 17248 11815
rect 20714 11812 20720 11824
rect 17190 11775 17248 11781
rect 19352 11784 20720 11812
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14608 11716 14657 11744
rect 14608 11704 14614 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11744 14887 11747
rect 15102 11744 15108 11756
rect 14875 11716 15108 11744
rect 14875 11713 14887 11716
rect 14829 11707 14887 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 17494 11744 17500 11756
rect 16163 11716 17500 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 5644 11648 6500 11676
rect 8205 11679 8263 11685
rect 5644 11617 5672 11648
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8294 11676 8300 11688
rect 8251 11648 8300 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11676 14151 11679
rect 14568 11676 14596 11704
rect 14139 11648 14596 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11577 5687 11611
rect 15488 11608 15516 11707
rect 15948 11676 15976 11707
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 19352 11753 19380 11784
rect 20714 11772 20720 11784
rect 20772 11812 20778 11824
rect 22278 11812 22284 11824
rect 20772 11784 22284 11812
rect 20772 11772 20778 11784
rect 22278 11772 22284 11784
rect 22336 11812 22342 11824
rect 25590 11812 25596 11824
rect 22336 11784 25596 11812
rect 22336 11772 22342 11784
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19604 11747 19662 11753
rect 19604 11713 19616 11747
rect 19650 11744 19662 11747
rect 20530 11744 20536 11756
rect 19650 11716 20536 11744
rect 19650 11713 19662 11716
rect 19604 11707 19662 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11744 22063 11747
rect 22094 11744 22100 11756
rect 22051 11716 22100 11744
rect 22051 11713 22063 11716
rect 22005 11707 22063 11713
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 22833 11707 22891 11713
rect 16666 11676 16672 11688
rect 15948 11648 16672 11676
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 16942 11676 16948 11688
rect 16816 11648 16948 11676
rect 16816 11636 16822 11648
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 21910 11636 21916 11688
rect 21968 11676 21974 11688
rect 22204 11676 22232 11707
rect 21968 11648 22232 11676
rect 22848 11676 22876 11707
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23658 11744 23664 11756
rect 23619 11716 23664 11744
rect 23658 11704 23664 11716
rect 23716 11704 23722 11756
rect 24412 11753 24440 11784
rect 25590 11772 25596 11784
rect 25648 11812 25654 11824
rect 26602 11812 26608 11824
rect 25648 11784 26608 11812
rect 25648 11772 25654 11784
rect 26602 11772 26608 11784
rect 26660 11772 26666 11824
rect 27522 11812 27528 11824
rect 26988 11784 27528 11812
rect 24670 11753 24676 11756
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 24664 11707 24676 11753
rect 24728 11744 24734 11756
rect 26418 11744 26424 11756
rect 24728 11716 24764 11744
rect 26379 11716 26424 11744
rect 24670 11704 24676 11707
rect 24728 11704 24734 11716
rect 26418 11704 26424 11716
rect 26476 11704 26482 11756
rect 26988 11753 27016 11784
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 29080 11815 29138 11821
rect 29080 11781 29092 11815
rect 29126 11812 29138 11815
rect 30558 11812 30564 11824
rect 29126 11784 30564 11812
rect 29126 11781 29138 11784
rect 29080 11775 29138 11781
rect 30558 11772 30564 11784
rect 30616 11772 30622 11824
rect 26973 11747 27031 11753
rect 26973 11713 26985 11747
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27062 11704 27068 11756
rect 27120 11744 27126 11756
rect 27229 11747 27287 11753
rect 27229 11744 27241 11747
rect 27120 11716 27241 11744
rect 27120 11704 27126 11716
rect 27229 11713 27241 11716
rect 27275 11713 27287 11747
rect 27540 11744 27568 11772
rect 30852 11753 30880 11852
rect 31018 11840 31024 11852
rect 31076 11840 31082 11892
rect 31662 11772 31668 11824
rect 31720 11812 31726 11824
rect 31720 11784 34928 11812
rect 31720 11772 31726 11784
rect 28813 11747 28871 11753
rect 28813 11744 28825 11747
rect 27540 11716 28825 11744
rect 27229 11707 27287 11713
rect 28813 11713 28825 11716
rect 28859 11713 28871 11747
rect 28813 11707 28871 11713
rect 30837 11747 30895 11753
rect 30837 11713 30849 11747
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 32766 11744 32772 11756
rect 32355 11716 32772 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 23750 11676 23756 11688
rect 22848 11648 23756 11676
rect 21968 11636 21974 11648
rect 23750 11636 23756 11648
rect 23808 11636 23814 11688
rect 16850 11608 16856 11620
rect 15488 11580 16856 11608
rect 5629 11571 5687 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 18598 11568 18604 11620
rect 18656 11608 18662 11620
rect 21818 11608 21824 11620
rect 18656 11580 19288 11608
rect 18656 11568 18662 11580
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6788 11512 7757 11540
rect 6788 11500 6794 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10376 11512 10517 11540
rect 10376 11500 10382 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13262 11540 13268 11552
rect 12943 11512 13268 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13357 11543 13415 11549
rect 13357 11509 13369 11543
rect 13403 11540 13415 11543
rect 14182 11540 14188 11552
rect 13403 11512 14188 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 14737 11543 14795 11549
rect 14737 11540 14749 11543
rect 14516 11512 14749 11540
rect 14516 11500 14522 11512
rect 14737 11509 14749 11512
rect 14783 11509 14795 11543
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 14737 11503 14795 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 18196 11512 18337 11540
rect 18196 11500 18202 11512
rect 18325 11509 18337 11512
rect 18371 11540 18383 11543
rect 19150 11540 19156 11552
rect 18371 11512 19156 11540
rect 18371 11509 18383 11512
rect 18325 11503 18383 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19260 11540 19288 11580
rect 20640 11580 21496 11608
rect 21731 11580 21824 11608
rect 20640 11540 20668 11580
rect 19260 11512 20668 11540
rect 20717 11543 20775 11549
rect 20717 11509 20729 11543
rect 20763 11540 20775 11543
rect 21358 11540 21364 11552
rect 20763 11512 21364 11540
rect 20763 11509 20775 11512
rect 20717 11503 20775 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21468 11540 21496 11580
rect 21818 11568 21824 11580
rect 21876 11608 21882 11620
rect 22002 11608 22008 11620
rect 21876 11580 22008 11608
rect 21876 11568 21882 11580
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 26878 11608 26884 11620
rect 22296 11580 23612 11608
rect 22296 11540 22324 11580
rect 21468 11512 22324 11540
rect 22554 11500 22560 11552
rect 22612 11540 22618 11552
rect 23477 11543 23535 11549
rect 23477 11540 23489 11543
rect 22612 11512 23489 11540
rect 22612 11500 22618 11512
rect 23477 11509 23489 11512
rect 23523 11509 23535 11543
rect 23584 11540 23612 11580
rect 25700 11580 26884 11608
rect 25700 11540 25728 11580
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 23584 11512 25728 11540
rect 23477 11503 23535 11509
rect 25774 11500 25780 11552
rect 25832 11540 25838 11552
rect 26234 11540 26240 11552
rect 25832 11512 25877 11540
rect 26195 11512 26240 11540
rect 25832 11500 25838 11512
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 28258 11500 28264 11552
rect 28316 11540 28322 11552
rect 28353 11543 28411 11549
rect 28353 11540 28365 11543
rect 28316 11512 28365 11540
rect 28316 11500 28322 11512
rect 28353 11509 28365 11512
rect 28399 11509 28411 11543
rect 28828 11540 28856 11707
rect 32766 11704 32772 11716
rect 32824 11704 32830 11756
rect 33060 11753 33088 11784
rect 34900 11753 34928 11784
rect 33045 11747 33103 11753
rect 33045 11713 33057 11747
rect 33091 11713 33103 11747
rect 33301 11747 33359 11753
rect 33301 11744 33313 11747
rect 33045 11707 33103 11713
rect 33152 11716 33313 11744
rect 30653 11679 30711 11685
rect 30653 11645 30665 11679
rect 30699 11676 30711 11679
rect 30926 11676 30932 11688
rect 30699 11648 30932 11676
rect 30699 11645 30711 11648
rect 30653 11639 30711 11645
rect 30926 11636 30932 11648
rect 30984 11636 30990 11688
rect 32585 11679 32643 11685
rect 32585 11645 32597 11679
rect 32631 11676 32643 11679
rect 32950 11676 32956 11688
rect 32631 11648 32956 11676
rect 32631 11645 32643 11648
rect 32585 11639 32643 11645
rect 32950 11636 32956 11648
rect 33008 11636 33014 11688
rect 33152 11676 33180 11716
rect 33301 11713 33313 11716
rect 33347 11713 33359 11747
rect 33301 11707 33359 11713
rect 34885 11747 34943 11753
rect 34885 11713 34897 11747
rect 34931 11713 34943 11747
rect 35141 11747 35199 11753
rect 35141 11744 35153 11747
rect 34885 11707 34943 11713
rect 34992 11716 35153 11744
rect 33060 11648 33180 11676
rect 31202 11608 31208 11620
rect 30116 11580 31208 11608
rect 29546 11540 29552 11552
rect 28828 11512 29552 11540
rect 28353 11503 28411 11509
rect 29546 11500 29552 11512
rect 29604 11540 29610 11552
rect 30116 11540 30144 11580
rect 31202 11568 31208 11580
rect 31260 11568 31266 11620
rect 32125 11611 32183 11617
rect 32125 11577 32137 11611
rect 32171 11608 32183 11611
rect 33060 11608 33088 11648
rect 34146 11636 34152 11688
rect 34204 11676 34210 11688
rect 34992 11676 35020 11716
rect 35141 11713 35153 11716
rect 35187 11713 35199 11747
rect 35141 11707 35199 11713
rect 34204 11648 35020 11676
rect 34204 11636 34210 11648
rect 32171 11580 33088 11608
rect 32171 11577 32183 11580
rect 32125 11571 32183 11577
rect 29604 11512 30144 11540
rect 32493 11543 32551 11549
rect 29604 11500 29610 11512
rect 32493 11509 32505 11543
rect 32539 11540 32551 11543
rect 33318 11540 33324 11552
rect 32539 11512 33324 11540
rect 32539 11509 32551 11512
rect 32493 11503 32551 11509
rect 33318 11500 33324 11512
rect 33376 11500 33382 11552
rect 34422 11540 34428 11552
rect 34383 11512 34428 11540
rect 34422 11500 34428 11512
rect 34480 11500 34486 11552
rect 36262 11540 36268 11552
rect 36223 11512 36268 11540
rect 36262 11500 36268 11512
rect 36320 11500 36326 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 7800 11308 8401 11336
rect 7800 11296 7806 11308
rect 8389 11305 8401 11308
rect 8435 11305 8447 11339
rect 8389 11299 8447 11305
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11336 12590 11348
rect 12710 11336 12716 11348
rect 12584 11308 12716 11336
rect 12584 11296 12590 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 14056 11308 14473 11336
rect 14056 11296 14062 11308
rect 14461 11305 14473 11308
rect 14507 11336 14519 11339
rect 15746 11336 15752 11348
rect 14507 11308 15752 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 16724 11308 18061 11336
rect 16724 11296 16730 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 18049 11299 18107 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 23658 11336 23664 11348
rect 22787 11308 23664 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24670 11336 24676 11348
rect 24631 11308 24676 11336
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 25038 11336 25044 11348
rect 24999 11308 25044 11336
rect 25038 11296 25044 11308
rect 25096 11336 25102 11348
rect 25866 11336 25872 11348
rect 25096 11308 25872 11336
rect 25096 11296 25102 11308
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 26973 11339 27031 11345
rect 26973 11305 26985 11339
rect 27019 11336 27031 11339
rect 27062 11336 27068 11348
rect 27019 11308 27068 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 27341 11339 27399 11345
rect 27341 11305 27353 11339
rect 27387 11336 27399 11339
rect 27706 11336 27712 11348
rect 27387 11308 27712 11336
rect 27387 11305 27399 11308
rect 27341 11299 27399 11305
rect 27706 11296 27712 11308
rect 27764 11296 27770 11348
rect 28626 11296 28632 11348
rect 28684 11336 28690 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 28684 11308 29929 11336
rect 28684 11296 28690 11308
rect 29917 11305 29929 11308
rect 29963 11305 29975 11339
rect 29917 11299 29975 11305
rect 30101 11339 30159 11345
rect 30101 11305 30113 11339
rect 30147 11336 30159 11339
rect 30742 11336 30748 11348
rect 30147 11308 30748 11336
rect 30147 11305 30159 11308
rect 30101 11299 30159 11305
rect 30742 11296 30748 11308
rect 30800 11296 30806 11348
rect 33965 11339 34023 11345
rect 33965 11305 33977 11339
rect 34011 11336 34023 11339
rect 34146 11336 34152 11348
rect 34011 11308 34152 11336
rect 34011 11305 34023 11308
rect 33965 11299 34023 11305
rect 34146 11296 34152 11308
rect 34204 11296 34210 11348
rect 14826 11268 14832 11280
rect 11440 11240 14832 11268
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9674 11200 9680 11212
rect 9171 11172 9680 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9646 11160 9680 11172
rect 9732 11160 9738 11212
rect 10410 11200 10416 11212
rect 10371 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 7024 11132 7052 11160
rect 5215 11104 7052 11132
rect 7276 11135 7334 11141
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 7276 11101 7288 11135
rect 7322 11132 7334 11135
rect 7650 11132 7656 11144
rect 7322 11104 7656 11132
rect 7322 11101 7334 11104
rect 7276 11095 7334 11101
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 9398 11132 9404 11144
rect 9359 11104 9404 11132
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9646 11132 9674 11160
rect 11440 11132 11468 11240
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 17313 11271 17371 11277
rect 17313 11237 17325 11271
rect 17359 11268 17371 11271
rect 18230 11268 18236 11280
rect 17359 11240 18236 11268
rect 17359 11237 17371 11240
rect 17313 11231 17371 11237
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 24302 11228 24308 11280
rect 24360 11268 24366 11280
rect 26329 11271 26387 11277
rect 26329 11268 26341 11271
rect 24360 11240 26341 11268
rect 24360 11228 24366 11240
rect 26329 11237 26341 11240
rect 26375 11237 26387 11271
rect 26329 11231 26387 11237
rect 26878 11228 26884 11280
rect 26936 11268 26942 11280
rect 33870 11268 33876 11280
rect 26936 11240 33876 11268
rect 26936 11228 26942 11240
rect 33870 11228 33876 11240
rect 33928 11228 33934 11280
rect 12618 11200 12624 11212
rect 12268 11172 12624 11200
rect 12268 11141 12296 11172
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13320 11172 14136 11200
rect 13320 11160 13326 11172
rect 14108 11141 14136 11172
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18414 11200 18420 11212
rect 18196 11172 18276 11200
rect 18375 11172 18420 11200
rect 18196 11160 18202 11172
rect 9646 11104 11468 11132
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14093 11095 14151 11101
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11132 15163 11135
rect 15372 11135 15430 11141
rect 15151 11104 15240 11132
rect 15151 11101 15163 11104
rect 15105 11095 15163 11101
rect 5436 11067 5494 11073
rect 5436 11033 5448 11067
rect 5482 11064 5494 11067
rect 5626 11064 5632 11076
rect 5482 11036 5632 11064
rect 5482 11033 5494 11036
rect 5436 11027 5494 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 10686 11073 10692 11076
rect 10680 11064 10692 11073
rect 10647 11036 10692 11064
rect 10680 11027 10692 11036
rect 10686 11024 10692 11027
rect 10744 11024 10750 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13357 11067 13415 11073
rect 13357 11064 13369 11067
rect 13228 11036 13369 11064
rect 13228 11024 13234 11036
rect 13357 11033 13369 11036
rect 13403 11033 13415 11067
rect 13357 11027 13415 11033
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 15212 11064 15240 11104
rect 15372 11101 15384 11135
rect 15418 11101 15430 11135
rect 15372 11095 15430 11101
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 18046 11132 18052 11144
rect 17635 11104 18052 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 13587 11036 15240 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11480 10968 11805 10996
rect 11480 10956 11486 10968
rect 11793 10965 11805 10968
rect 11839 10965 11851 10999
rect 11793 10959 11851 10965
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 13556 10996 13584 11027
rect 14642 10996 14648 11008
rect 12400 10968 13584 10996
rect 14603 10968 14648 10996
rect 12400 10956 12406 10968
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15212 10996 15240 11036
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15396 11064 15424 11095
rect 18046 11092 18052 11104
rect 18104 11132 18110 11144
rect 18248 11141 18276 11172
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 22370 11200 22376 11212
rect 20036 11172 22376 11200
rect 20036 11160 20042 11172
rect 18233 11135 18291 11141
rect 18104 11104 18184 11132
rect 18104 11092 18110 11104
rect 16758 11064 16764 11076
rect 15344 11036 15424 11064
rect 15488 11036 16764 11064
rect 15344 11024 15350 11036
rect 15488 10996 15516 11036
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 17954 11064 17960 11076
rect 17359 11036 17960 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18156 11064 18184 11104
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18509 11135 18567 11141
rect 18380 11104 18425 11132
rect 18380 11092 18386 11104
rect 18509 11101 18521 11135
rect 18555 11132 18567 11135
rect 18598 11132 18604 11144
rect 18555 11104 18604 11132
rect 18555 11101 18567 11104
rect 18509 11095 18567 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19426 11132 19432 11144
rect 19291 11104 19432 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11132 20775 11135
rect 20806 11132 20812 11144
rect 20763 11104 20812 11132
rect 20763 11101 20775 11104
rect 20717 11095 20775 11101
rect 18340 11064 18368 11092
rect 19536 11064 19564 11095
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 21192 11141 21220 11172
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 25665 11203 25723 11209
rect 25665 11200 25677 11203
rect 24872 11172 25677 11200
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 22186 11132 22192 11144
rect 21407 11104 22192 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 23014 11132 23020 11144
rect 22388 11104 23020 11132
rect 18156 11036 19564 11064
rect 20898 11024 20904 11076
rect 20956 11064 20962 11076
rect 22388 11073 22416 11104
rect 23014 11092 23020 11104
rect 23072 11132 23078 11144
rect 24872 11141 24900 11172
rect 25665 11169 25677 11172
rect 25711 11169 25723 11203
rect 25665 11163 25723 11169
rect 26142 11160 26148 11212
rect 26200 11200 26206 11212
rect 27433 11203 27491 11209
rect 26200 11172 26648 11200
rect 26200 11160 26206 11172
rect 23385 11135 23443 11141
rect 23385 11132 23397 11135
rect 23072 11104 23397 11132
rect 23072 11092 23078 11104
rect 23385 11101 23397 11104
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 25130 11132 25136 11144
rect 25091 11104 25136 11132
rect 24857 11095 24915 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25240 11104 25820 11132
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20956 11036 21281 11064
rect 20956 11024 20962 11036
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21269 11027 21327 11033
rect 22373 11067 22431 11073
rect 22373 11033 22385 11067
rect 22419 11033 22431 11067
rect 22373 11027 22431 11033
rect 22557 11067 22615 11073
rect 22557 11033 22569 11067
rect 22603 11064 22615 11067
rect 23198 11064 23204 11076
rect 22603 11036 23204 11064
rect 22603 11033 22615 11036
rect 22557 11027 22615 11033
rect 23198 11024 23204 11036
rect 23256 11024 23262 11076
rect 23569 11067 23627 11073
rect 23569 11033 23581 11067
rect 23615 11064 23627 11067
rect 23753 11067 23811 11073
rect 23615 11036 23704 11064
rect 23615 11033 23627 11036
rect 23569 11027 23627 11033
rect 16482 10996 16488 11008
rect 15212 10968 15516 10996
rect 16443 10968 16488 10996
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 17497 10999 17555 11005
rect 17497 10965 17509 10999
rect 17543 10996 17555 10999
rect 17678 10996 17684 11008
rect 17543 10968 17684 10996
rect 17543 10965 17555 10968
rect 17497 10959 17555 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 23676 10996 23704 11036
rect 23753 11033 23765 11067
rect 23799 11064 23811 11067
rect 25240 11064 25268 11104
rect 23799 11036 25268 11064
rect 23799 11033 23811 11036
rect 23753 11027 23811 11033
rect 25314 11024 25320 11076
rect 25372 11064 25378 11076
rect 25593 11067 25651 11073
rect 25372 11036 25544 11064
rect 25372 11024 25378 11036
rect 25038 10996 25044 11008
rect 23676 10968 25044 10996
rect 25038 10956 25044 10968
rect 25096 10956 25102 11008
rect 25516 10996 25544 11036
rect 25593 11033 25605 11067
rect 25639 11064 25651 11067
rect 25682 11064 25688 11076
rect 25639 11036 25688 11064
rect 25639 11033 25651 11036
rect 25593 11027 25651 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 25792 11064 25820 11104
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 26513 11135 26571 11141
rect 25924 11104 25969 11132
rect 25924 11092 25930 11104
rect 26513 11101 26525 11135
rect 26559 11101 26571 11135
rect 26513 11095 26571 11101
rect 26528 11064 26556 11095
rect 25792 11036 26556 11064
rect 26620 11064 26648 11172
rect 27433 11169 27445 11203
rect 27479 11200 27491 11203
rect 28258 11200 28264 11212
rect 27479 11172 28264 11200
rect 27479 11169 27491 11172
rect 27433 11163 27491 11169
rect 28258 11160 28264 11172
rect 28316 11160 28322 11212
rect 29549 11203 29607 11209
rect 29549 11169 29561 11203
rect 29595 11200 29607 11203
rect 29914 11200 29920 11212
rect 29595 11172 29920 11200
rect 29595 11169 29607 11172
rect 29549 11163 29607 11169
rect 29914 11160 29920 11172
rect 29972 11160 29978 11212
rect 30929 11203 30987 11209
rect 30929 11200 30941 11203
rect 30024 11172 30941 11200
rect 27154 11132 27160 11144
rect 27115 11104 27160 11132
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 27338 11092 27344 11144
rect 27396 11132 27402 11144
rect 28077 11135 28135 11141
rect 28077 11132 28089 11135
rect 27396 11104 28089 11132
rect 27396 11092 27402 11104
rect 28077 11101 28089 11104
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11132 28779 11135
rect 28902 11132 28908 11144
rect 28767 11104 28908 11132
rect 28767 11101 28779 11104
rect 28721 11095 28779 11101
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 28997 11135 29055 11141
rect 28997 11101 29009 11135
rect 29043 11132 29055 11135
rect 29822 11132 29828 11144
rect 29043 11104 29828 11132
rect 29043 11101 29055 11104
rect 28997 11095 29055 11101
rect 29822 11092 29828 11104
rect 29880 11132 29886 11144
rect 30024 11132 30052 11172
rect 30929 11169 30941 11172
rect 30975 11169 30987 11203
rect 32674 11200 32680 11212
rect 32635 11172 32680 11200
rect 30929 11163 30987 11169
rect 32674 11160 32680 11172
rect 32732 11160 32738 11212
rect 29880 11104 30052 11132
rect 29880 11092 29886 11104
rect 30650 11092 30656 11144
rect 30708 11132 30714 11144
rect 30745 11135 30803 11141
rect 30745 11132 30757 11135
rect 30708 11104 30757 11132
rect 30708 11092 30714 11104
rect 30745 11101 30757 11104
rect 30791 11101 30803 11135
rect 31018 11132 31024 11144
rect 30745 11095 30803 11101
rect 30852 11104 31024 11132
rect 28537 11067 28595 11073
rect 26620 11036 27936 11064
rect 25774 10996 25780 11008
rect 25516 10968 25780 10996
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 25866 10956 25872 11008
rect 25924 10996 25930 11008
rect 27338 10996 27344 11008
rect 25924 10968 27344 10996
rect 25924 10956 25930 10968
rect 27338 10956 27344 10968
rect 27396 10956 27402 11008
rect 27908 11005 27936 11036
rect 28537 11033 28549 11067
rect 28583 11064 28595 11067
rect 29917 11067 29975 11073
rect 29917 11064 29929 11067
rect 28583 11036 29929 11064
rect 28583 11033 28595 11036
rect 28537 11027 28595 11033
rect 29917 11033 29929 11036
rect 29963 11033 29975 11067
rect 30852 11064 30880 11104
rect 31018 11092 31024 11104
rect 31076 11132 31082 11144
rect 31757 11135 31815 11141
rect 31757 11132 31769 11135
rect 31076 11104 31769 11132
rect 31076 11092 31082 11104
rect 31757 11101 31769 11104
rect 31803 11101 31815 11135
rect 31757 11095 31815 11101
rect 32953 11135 33011 11141
rect 32953 11101 32965 11135
rect 32999 11132 33011 11135
rect 33502 11132 33508 11144
rect 32999 11104 33508 11132
rect 32999 11101 33011 11104
rect 32953 11095 33011 11101
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 33962 11132 33968 11144
rect 33923 11104 33968 11132
rect 33962 11092 33968 11104
rect 34020 11092 34026 11144
rect 34146 11132 34152 11144
rect 34107 11104 34152 11132
rect 34146 11092 34152 11104
rect 34204 11092 34210 11144
rect 31573 11067 31631 11073
rect 31573 11064 31585 11067
rect 29917 11027 29975 11033
rect 30392 11036 30880 11064
rect 30944 11036 31585 11064
rect 27893 10999 27951 11005
rect 27893 10965 27905 10999
rect 27939 10965 27951 10999
rect 27893 10959 27951 10965
rect 28905 10999 28963 11005
rect 28905 10965 28917 10999
rect 28951 10996 28963 10999
rect 30392 10996 30420 11036
rect 30944 11008 30972 11036
rect 31573 11033 31585 11036
rect 31619 11033 31631 11067
rect 31573 11027 31631 11033
rect 30558 10996 30564 11008
rect 28951 10968 30420 10996
rect 30519 10968 30564 10996
rect 28951 10965 28963 10968
rect 28905 10959 28963 10965
rect 30558 10956 30564 10968
rect 30616 10956 30622 11008
rect 30926 10956 30932 11008
rect 30984 10956 30990 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 5626 10792 5632 10804
rect 5587 10764 5632 10792
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 6972 10764 7297 10792
rect 6972 10752 6978 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9582 10792 9588 10804
rect 8352 10764 9588 10792
rect 8352 10752 8358 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9950 10792 9956 10804
rect 9911 10764 9956 10792
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11330 10792 11336 10804
rect 11011 10764 11336 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 13725 10795 13783 10801
rect 11900 10764 13676 10792
rect 8113 10727 8171 10733
rect 8113 10724 8125 10727
rect 5828 10696 8125 10724
rect 5828 10665 5856 10696
rect 8113 10693 8125 10696
rect 8159 10693 8171 10727
rect 10318 10724 10324 10736
rect 8113 10687 8171 10693
rect 8588 10696 10324 10724
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 5813 10619 5871 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7190 10656 7196 10668
rect 7147 10628 7196 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 7024 10588 7052 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 7926 10656 7932 10668
rect 7887 10628 7932 10656
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8588 10665 8616 10696
rect 10318 10684 10324 10696
rect 10376 10724 10382 10736
rect 11900 10733 11928 10764
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 10376 10696 11713 10724
rect 10376 10684 10382 10696
rect 11701 10693 11713 10696
rect 11747 10693 11759 10727
rect 11701 10687 11759 10693
rect 11885 10727 11943 10733
rect 11885 10693 11897 10727
rect 11931 10693 11943 10727
rect 11885 10687 11943 10693
rect 12434 10684 12440 10736
rect 12492 10724 12498 10736
rect 12590 10727 12648 10733
rect 12590 10724 12602 10727
rect 12492 10696 12602 10724
rect 12492 10684 12498 10696
rect 12590 10693 12602 10696
rect 12636 10693 12648 10727
rect 12590 10687 12648 10693
rect 12710 10684 12716 10736
rect 12768 10684 12774 10736
rect 13648 10724 13676 10764
rect 13725 10761 13737 10795
rect 13771 10792 13783 10795
rect 17678 10792 17684 10804
rect 13771 10764 14228 10792
rect 17591 10764 17684 10792
rect 13771 10761 13783 10764
rect 13725 10755 13783 10761
rect 13998 10724 14004 10736
rect 13648 10696 14004 10724
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8754 10656 8760 10668
rect 8715 10628 8760 10656
rect 8573 10619 8631 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9306 10656 9312 10668
rect 8987 10628 9312 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 2464 10560 7052 10588
rect 7745 10591 7803 10597
rect 2464 10548 2470 10560
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8294 10588 8300 10600
rect 7791 10560 8300 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 8864 10520 8892 10619
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 9769 10619 9827 10625
rect 9582 10588 9588 10600
rect 9543 10560 9588 10588
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 3292 10492 8892 10520
rect 9125 10523 9183 10529
rect 3292 10480 3298 10492
rect 9125 10489 9137 10523
rect 9171 10520 9183 10523
rect 9784 10520 9812 10619
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10796 10588 10824 10619
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11480 10628 11529 10656
rect 11480 10616 11486 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 12342 10656 12348 10668
rect 12303 10628 12348 10656
rect 11517 10619 11575 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12728 10656 12756 10684
rect 14200 10665 14228 10764
rect 17678 10752 17684 10764
rect 17736 10792 17742 10804
rect 18506 10792 18512 10804
rect 17736 10764 18512 10792
rect 17736 10752 17742 10764
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18969 10795 19027 10801
rect 18969 10761 18981 10795
rect 19015 10792 19027 10795
rect 19242 10792 19248 10804
rect 19015 10764 19248 10792
rect 19015 10761 19027 10764
rect 18969 10755 19027 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 22830 10792 22836 10804
rect 22664 10764 22836 10792
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 17402 10724 17408 10736
rect 14884 10696 17408 10724
rect 14884 10684 14890 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 18138 10724 18144 10736
rect 17543 10696 18144 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 18325 10727 18383 10733
rect 18325 10693 18337 10727
rect 18371 10724 18383 10727
rect 18414 10724 18420 10736
rect 18371 10696 18420 10724
rect 18371 10693 18383 10696
rect 18325 10687 18383 10693
rect 18414 10684 18420 10696
rect 18472 10724 18478 10736
rect 21358 10724 21364 10736
rect 18472 10696 19380 10724
rect 18472 10684 18478 10696
rect 12452 10628 12756 10656
rect 14185 10659 14243 10665
rect 12452 10588 12480 10628
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14366 10656 14372 10668
rect 14231 10628 14372 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 14424 10628 15485 10656
rect 14424 10616 14430 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15746 10656 15752 10668
rect 15707 10628 15752 10656
rect 15473 10619 15531 10625
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16040 10628 16681 10656
rect 10796 10560 12480 10588
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 14332 10560 14473 10588
rect 14332 10548 14338 10560
rect 14461 10557 14473 10560
rect 14507 10588 14519 10591
rect 15102 10588 15108 10600
rect 14507 10560 15108 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 15933 10591 15991 10597
rect 15933 10588 15945 10591
rect 15896 10560 15945 10588
rect 15896 10548 15902 10560
rect 15933 10557 15945 10560
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 9171 10492 9812 10520
rect 15120 10520 15148 10548
rect 16040 10520 16068 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 16942 10656 16948 10668
rect 16899 10628 16948 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10656 17831 10659
rect 18046 10656 18052 10668
rect 17819 10628 18052 10656
rect 17819 10625 17831 10628
rect 17773 10619 17831 10625
rect 18046 10616 18052 10628
rect 18104 10656 18110 10668
rect 19352 10665 19380 10696
rect 19444 10696 21364 10724
rect 19444 10665 19472 10696
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 21450 10684 21456 10736
rect 21508 10724 21514 10736
rect 22664 10733 22692 10764
rect 22830 10752 22836 10764
rect 22888 10792 22894 10804
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 22888 10764 25697 10792
rect 22888 10752 22894 10764
rect 25685 10761 25697 10764
rect 25731 10761 25743 10795
rect 28350 10792 28356 10804
rect 25685 10755 25743 10761
rect 26252 10764 28356 10792
rect 22649 10727 22707 10733
rect 21508 10696 22048 10724
rect 21508 10684 21514 10696
rect 19245 10659 19303 10665
rect 19245 10656 19257 10659
rect 18104 10628 19257 10656
rect 18104 10616 18110 10628
rect 19245 10625 19257 10628
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 19337 10659 19395 10665
rect 19337 10625 19349 10659
rect 19383 10625 19395 10659
rect 19337 10619 19395 10625
rect 19429 10659 19487 10665
rect 19429 10625 19441 10659
rect 19475 10625 19487 10659
rect 21174 10656 21180 10668
rect 21135 10628 21180 10656
rect 19429 10619 19487 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 21818 10656 21824 10668
rect 21779 10628 21824 10656
rect 21818 10616 21824 10628
rect 21876 10616 21882 10668
rect 22020 10665 22048 10696
rect 22649 10693 22661 10727
rect 22695 10693 22707 10727
rect 22649 10687 22707 10693
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10724 22799 10727
rect 23566 10724 23572 10736
rect 22787 10696 23572 10724
rect 22787 10693 22799 10696
rect 22741 10687 22799 10693
rect 23566 10684 23572 10696
rect 23624 10684 23630 10736
rect 23934 10724 23940 10736
rect 23676 10696 23940 10724
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22152 10628 22477 10656
rect 22152 10616 22158 10628
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10656 22891 10659
rect 23106 10656 23112 10668
rect 22879 10628 23112 10656
rect 22879 10625 22891 10628
rect 22833 10619 22891 10625
rect 23106 10616 23112 10628
rect 23164 10616 23170 10668
rect 23676 10665 23704 10696
rect 23934 10684 23940 10696
rect 23992 10684 23998 10736
rect 23661 10659 23719 10665
rect 23661 10625 23673 10659
rect 23707 10625 23719 10659
rect 23842 10656 23848 10668
rect 23803 10628 23848 10656
rect 23661 10619 23719 10625
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 24857 10659 24915 10665
rect 24857 10656 24869 10659
rect 24728 10628 24869 10656
rect 24728 10616 24734 10628
rect 24857 10625 24869 10628
rect 24903 10625 24915 10659
rect 25590 10656 25596 10668
rect 25551 10628 25596 10656
rect 24857 10619 24915 10625
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 26252 10665 26280 10764
rect 28350 10752 28356 10764
rect 28408 10792 28414 10804
rect 30926 10792 30932 10804
rect 28408 10764 30820 10792
rect 30887 10764 30932 10792
rect 28408 10752 28414 10764
rect 28442 10724 28448 10736
rect 26344 10696 28448 10724
rect 26237 10659 26295 10665
rect 26237 10625 26249 10659
rect 26283 10625 26295 10659
rect 26237 10619 26295 10625
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16163 10560 19104 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 17494 10520 17500 10532
rect 15120 10492 16068 10520
rect 16132 10492 16988 10520
rect 17455 10492 17500 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 9490 10452 9496 10464
rect 2924 10424 9496 10452
rect 2924 10412 2930 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 16132 10452 16160 10492
rect 16960 10464 16988 10492
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 18506 10520 18512 10532
rect 18467 10492 18512 10520
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 19076 10520 19104 10560
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19208 10560 19253 10588
rect 19306 10560 19472 10588
rect 19208 10548 19214 10560
rect 19306 10520 19334 10560
rect 19076 10492 19334 10520
rect 19444 10520 19472 10560
rect 19886 10548 19892 10600
rect 19944 10588 19950 10600
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19944 10560 19993 10588
rect 19944 10548 19950 10560
rect 19981 10557 19993 10560
rect 20027 10588 20039 10591
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 20027 10560 23949 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 20346 10520 20352 10532
rect 19444 10492 20352 10520
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 20993 10523 21051 10529
rect 20993 10489 21005 10523
rect 21039 10520 21051 10523
rect 22462 10520 22468 10532
rect 21039 10492 22468 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 24210 10480 24216 10532
rect 24268 10520 24274 10532
rect 26237 10523 26295 10529
rect 26237 10520 26249 10523
rect 24268 10492 26249 10520
rect 24268 10480 24274 10492
rect 26237 10489 26249 10492
rect 26283 10489 26295 10523
rect 26237 10483 26295 10489
rect 15436 10424 16160 10452
rect 15436 10412 15442 10424
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16632 10424 16773 10452
rect 16632 10412 16638 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 19886 10452 19892 10464
rect 17000 10424 19892 10452
rect 17000 10412 17006 10424
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 21821 10455 21879 10461
rect 21821 10421 21833 10455
rect 21867 10452 21879 10455
rect 22922 10452 22928 10464
rect 21867 10424 22928 10452
rect 21867 10421 21879 10424
rect 21821 10415 21879 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23017 10455 23075 10461
rect 23017 10421 23029 10455
rect 23063 10452 23075 10455
rect 23198 10452 23204 10464
rect 23063 10424 23204 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 23474 10452 23480 10464
rect 23435 10424 23480 10452
rect 23474 10412 23480 10424
rect 23532 10412 23538 10464
rect 24949 10455 25007 10461
rect 24949 10421 24961 10455
rect 24995 10452 25007 10455
rect 25498 10452 25504 10464
rect 24995 10424 25504 10452
rect 24995 10421 25007 10424
rect 24949 10415 25007 10421
rect 25498 10412 25504 10424
rect 25556 10412 25562 10464
rect 25682 10412 25688 10464
rect 25740 10452 25746 10464
rect 26344 10452 26372 10696
rect 28442 10684 28448 10696
rect 28500 10684 28506 10736
rect 29816 10727 29874 10733
rect 29816 10693 29828 10727
rect 29862 10724 29874 10727
rect 30558 10724 30564 10736
rect 29862 10696 30564 10724
rect 29862 10693 29874 10696
rect 29816 10687 29874 10693
rect 30558 10684 30564 10696
rect 30616 10684 30622 10736
rect 30792 10724 30820 10764
rect 30926 10752 30932 10764
rect 30984 10752 30990 10804
rect 32953 10795 33011 10801
rect 32953 10761 32965 10795
rect 32999 10792 33011 10795
rect 33134 10792 33140 10804
rect 32999 10764 33140 10792
rect 32999 10761 33011 10764
rect 32953 10755 33011 10761
rect 33134 10752 33140 10764
rect 33192 10792 33198 10804
rect 33689 10795 33747 10801
rect 33689 10792 33701 10795
rect 33192 10764 33701 10792
rect 33192 10752 33198 10764
rect 33689 10761 33701 10764
rect 33735 10792 33747 10795
rect 34238 10792 34244 10804
rect 33735 10764 34244 10792
rect 33735 10761 33747 10764
rect 33689 10755 33747 10761
rect 34238 10752 34244 10764
rect 34296 10792 34302 10804
rect 34296 10764 34560 10792
rect 34296 10752 34302 10764
rect 31386 10724 31392 10736
rect 30792 10696 31392 10724
rect 31386 10684 31392 10696
rect 31444 10684 31450 10736
rect 33318 10724 33324 10736
rect 33060 10696 33324 10724
rect 26421 10659 26479 10665
rect 26421 10625 26433 10659
rect 26467 10656 26479 10659
rect 26510 10656 26516 10668
rect 26467 10628 26516 10656
rect 26467 10625 26479 10628
rect 26421 10619 26479 10625
rect 26510 10616 26516 10628
rect 26568 10616 26574 10668
rect 27065 10659 27123 10665
rect 27065 10625 27077 10659
rect 27111 10625 27123 10659
rect 27065 10619 27123 10625
rect 28169 10659 28227 10665
rect 28169 10625 28181 10659
rect 28215 10625 28227 10659
rect 28902 10656 28908 10668
rect 28863 10628 28908 10656
rect 28169 10619 28227 10625
rect 27080 10520 27108 10619
rect 28184 10588 28212 10619
rect 28902 10616 28908 10628
rect 28960 10616 28966 10668
rect 29546 10656 29552 10668
rect 29507 10628 29552 10656
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 29638 10616 29644 10668
rect 29696 10656 29702 10668
rect 29696 10628 30604 10656
rect 29696 10616 29702 10628
rect 30576 10588 30604 10628
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 31573 10659 31631 10665
rect 31573 10656 31585 10659
rect 30984 10628 31585 10656
rect 30984 10616 30990 10628
rect 31573 10625 31585 10628
rect 31619 10625 31631 10659
rect 31573 10619 31631 10625
rect 31662 10616 31668 10668
rect 31720 10656 31726 10668
rect 33060 10665 33088 10696
rect 33318 10684 33324 10696
rect 33376 10724 33382 10736
rect 33376 10696 33824 10724
rect 33376 10684 33382 10696
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 31720 10628 32321 10656
rect 31720 10616 31726 10628
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32769 10659 32827 10665
rect 32769 10625 32781 10659
rect 32815 10625 32827 10659
rect 32769 10619 32827 10625
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10625 33103 10659
rect 33410 10656 33416 10668
rect 33323 10628 33416 10656
rect 33045 10619 33103 10625
rect 32784 10588 32812 10619
rect 33336 10600 33364 10628
rect 33410 10616 33416 10628
rect 33468 10656 33474 10668
rect 33796 10665 33824 10696
rect 33505 10659 33563 10665
rect 33505 10656 33517 10659
rect 33468 10628 33517 10656
rect 33468 10616 33474 10628
rect 33505 10625 33517 10628
rect 33551 10625 33563 10659
rect 33505 10619 33563 10625
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 33781 10619 33839 10625
rect 34241 10659 34299 10665
rect 34241 10625 34253 10659
rect 34287 10656 34299 10659
rect 34422 10656 34428 10668
rect 34287 10628 34428 10656
rect 34287 10625 34299 10628
rect 34241 10619 34299 10625
rect 34422 10616 34428 10628
rect 34480 10616 34486 10668
rect 34532 10665 34560 10764
rect 34517 10659 34575 10665
rect 34517 10625 34529 10659
rect 34563 10625 34575 10659
rect 34517 10619 34575 10625
rect 35713 10659 35771 10665
rect 35713 10625 35725 10659
rect 35759 10625 35771 10659
rect 35713 10619 35771 10625
rect 28184 10560 29132 10588
rect 30576 10560 32812 10588
rect 29104 10532 29132 10560
rect 33318 10548 33324 10600
rect 33376 10548 33382 10600
rect 29086 10520 29092 10532
rect 27080 10492 28304 10520
rect 29047 10492 29092 10520
rect 25740 10424 26372 10452
rect 25740 10412 25746 10424
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 28276 10461 28304 10492
rect 29086 10480 29092 10492
rect 29144 10480 29150 10532
rect 30558 10480 30564 10532
rect 30616 10520 30622 10532
rect 32766 10520 32772 10532
rect 30616 10492 32628 10520
rect 32727 10492 32772 10520
rect 30616 10480 30622 10492
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 26660 10424 27169 10452
rect 26660 10412 26666 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27157 10415 27215 10421
rect 28261 10455 28319 10461
rect 28261 10421 28273 10455
rect 28307 10452 28319 10455
rect 30742 10452 30748 10464
rect 28307 10424 30748 10452
rect 28307 10421 28319 10424
rect 28261 10415 28319 10421
rect 30742 10412 30748 10424
rect 30800 10412 30806 10464
rect 30834 10412 30840 10464
rect 30892 10452 30898 10464
rect 31389 10455 31447 10461
rect 31389 10452 31401 10455
rect 30892 10424 31401 10452
rect 30892 10412 30898 10424
rect 31389 10421 31401 10424
rect 31435 10421 31447 10455
rect 31389 10415 31447 10421
rect 31938 10412 31944 10464
rect 31996 10452 32002 10464
rect 32125 10455 32183 10461
rect 32125 10452 32137 10455
rect 31996 10424 32137 10452
rect 31996 10412 32002 10424
rect 32125 10421 32137 10424
rect 32171 10421 32183 10455
rect 32600 10452 32628 10492
rect 32766 10480 32772 10492
rect 32824 10480 32830 10532
rect 33505 10523 33563 10529
rect 33505 10489 33517 10523
rect 33551 10520 33563 10523
rect 34146 10520 34152 10532
rect 33551 10492 34152 10520
rect 33551 10489 33563 10492
rect 33505 10483 33563 10489
rect 34146 10480 34152 10492
rect 34204 10480 34210 10532
rect 35728 10520 35756 10619
rect 34256 10492 35756 10520
rect 34256 10452 34284 10492
rect 32600 10424 34284 10452
rect 32125 10415 32183 10421
rect 34606 10412 34612 10464
rect 34664 10452 34670 10464
rect 35529 10455 35587 10461
rect 35529 10452 35541 10455
rect 34664 10424 35541 10452
rect 34664 10412 34670 10424
rect 35529 10421 35541 10424
rect 35575 10421 35587 10455
rect 35529 10415 35587 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7926 10248 7932 10260
rect 7147 10220 7932 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 8386 10248 8392 10260
rect 8251 10220 8392 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9766 10248 9772 10260
rect 9539 10220 9772 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11241 10251 11299 10257
rect 11241 10248 11253 10251
rect 11112 10220 11253 10248
rect 11112 10208 11118 10220
rect 11241 10217 11253 10220
rect 11287 10248 11299 10251
rect 12158 10248 12164 10260
rect 11287 10220 12164 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 13357 10251 13415 10257
rect 13357 10217 13369 10251
rect 13403 10248 13415 10251
rect 15378 10248 15384 10260
rect 13403 10220 15384 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 4764 10152 7052 10180
rect 4764 10140 4770 10152
rect 7024 10112 7052 10152
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 10321 10183 10379 10189
rect 7248 10152 8064 10180
rect 7248 10140 7254 10152
rect 7024 10084 7972 10112
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 6178 10044 6184 10056
rect 5307 10016 6184 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6656 10016 6837 10044
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5408 9948 5457 9976
rect 5408 9936 5414 9948
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6656 9976 6684 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7190 10044 7196 10056
rect 6963 10016 7196 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 7742 10044 7748 10056
rect 7699 10016 7748 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 7944 10053 7972 10084
rect 8036 10053 8064 10152
rect 10321 10149 10333 10183
rect 10367 10180 10379 10183
rect 10502 10180 10508 10192
rect 10367 10152 10508 10180
rect 10367 10149 10379 10152
rect 10321 10143 10379 10149
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 13372 10180 13400 10211
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18598 10248 18604 10260
rect 18012 10220 18604 10248
rect 18012 10208 18018 10220
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 21232 10220 22937 10248
rect 21232 10208 21238 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 28902 10248 28908 10260
rect 22925 10211 22983 10217
rect 25516 10220 28908 10248
rect 18322 10180 18328 10192
rect 10612 10152 13400 10180
rect 14476 10152 18328 10180
rect 10612 10112 10640 10152
rect 8956 10084 10640 10112
rect 8956 10053 8984 10084
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 9306 10044 9312 10056
rect 8941 10007 8999 10013
rect 9048 10016 9312 10044
rect 5868 9948 6684 9976
rect 6733 9979 6791 9985
rect 5868 9936 5874 9948
rect 6733 9945 6745 9979
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 7837 9979 7895 9985
rect 7837 9945 7849 9979
rect 7883 9945 7895 9979
rect 8036 9976 8064 10007
rect 9048 9976 9076 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11057 10007 11115 10013
rect 8036 9948 9076 9976
rect 9125 9979 9183 9985
rect 7837 9939 7895 9945
rect 9125 9945 9137 9979
rect 9171 9945 9183 9979
rect 9125 9939 9183 9945
rect 9217 9979 9275 9985
rect 9217 9945 9229 9979
rect 9263 9976 9275 9979
rect 9490 9976 9496 9988
rect 9263 9948 9496 9976
rect 9263 9945 9275 9948
rect 9217 9939 9275 9945
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 6362 9908 6368 9920
rect 5675 9880 6368 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6748 9908 6776 9939
rect 6914 9908 6920 9920
rect 6748 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9908 6978 9920
rect 7852 9908 7880 9939
rect 8754 9908 8760 9920
rect 6972 9880 8760 9908
rect 6972 9868 6978 9880
rect 8754 9868 8760 9880
rect 8812 9908 8818 9920
rect 9140 9908 9168 9939
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 10134 9976 10140 9988
rect 10095 9948 10140 9976
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 11072 9976 11100 10007
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 11974 10044 11980 10056
rect 11931 10016 11980 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 13262 10044 13268 10056
rect 13223 10016 13268 10044
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14476 10053 14504 10152
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 18782 10140 18788 10192
rect 18840 10180 18846 10192
rect 21637 10183 21695 10189
rect 21637 10180 21649 10183
rect 18840 10152 21649 10180
rect 18840 10140 18846 10152
rect 21637 10149 21649 10152
rect 21683 10180 21695 10183
rect 25516 10180 25544 10220
rect 28902 10208 28908 10220
rect 28960 10208 28966 10260
rect 29917 10251 29975 10257
rect 29917 10217 29929 10251
rect 29963 10248 29975 10251
rect 30650 10248 30656 10260
rect 29963 10220 30656 10248
rect 29963 10217 29975 10220
rect 29917 10211 29975 10217
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 31386 10208 31392 10260
rect 31444 10248 31450 10260
rect 32950 10248 32956 10260
rect 31444 10220 32956 10248
rect 31444 10208 31450 10220
rect 32950 10208 32956 10220
rect 33008 10208 33014 10260
rect 33410 10208 33416 10260
rect 33468 10248 33474 10260
rect 35989 10251 36047 10257
rect 35989 10248 36001 10251
rect 33468 10220 36001 10248
rect 33468 10208 33474 10220
rect 35989 10217 36001 10220
rect 36035 10217 36047 10251
rect 35989 10211 36047 10217
rect 21683 10152 25544 10180
rect 25869 10183 25927 10189
rect 21683 10149 21695 10152
rect 21637 10143 21695 10149
rect 25869 10149 25881 10183
rect 25915 10149 25927 10183
rect 28442 10180 28448 10192
rect 28403 10152 28448 10180
rect 25869 10143 25927 10149
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 25590 10112 25596 10124
rect 15068 10084 20392 10112
rect 15068 10072 15074 10084
rect 14461 10047 14519 10053
rect 14240 10016 14412 10044
rect 14240 10004 14246 10016
rect 14274 9976 14280 9988
rect 11072 9948 14280 9976
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14384 9976 14412 10016
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 14608 10016 14657 10044
rect 14608 10004 14614 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14826 10044 14832 10056
rect 14787 10016 14832 10044
rect 14645 10007 14703 10013
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15488 10016 15761 10044
rect 14384 9948 14596 9976
rect 8812 9880 9168 9908
rect 10781 9911 10839 9917
rect 8812 9868 8818 9880
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 11514 9908 11520 9920
rect 10827 9880 11520 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 14568 9917 14596 9948
rect 15102 9936 15108 9988
rect 15160 9976 15166 9988
rect 15488 9976 15516 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15896 10016 15945 10044
rect 15896 10004 15902 10016
rect 15933 10013 15945 10016
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 16390 10004 16396 10056
rect 16448 10044 16454 10056
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 16448 10016 16497 10044
rect 16448 10004 16454 10016
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16666 10044 16672 10056
rect 16627 10016 16672 10044
rect 16485 10007 16543 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17420 10016 18092 10044
rect 17420 9976 17448 10016
rect 15160 9948 15516 9976
rect 15580 9948 17448 9976
rect 17497 9979 17555 9985
rect 15160 9936 15166 9948
rect 15580 9917 15608 9948
rect 17497 9945 17509 9979
rect 17543 9976 17555 9979
rect 17954 9976 17960 9988
rect 17543 9948 17960 9976
rect 17543 9945 17555 9948
rect 17497 9939 17555 9945
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 11664 9880 12081 9908
rect 11664 9868 11670 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9877 14611 9911
rect 14553 9871 14611 9877
rect 15565 9911 15623 9917
rect 15565 9877 15577 9911
rect 15611 9877 15623 9911
rect 15565 9871 15623 9877
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 17512 9908 17540 9939
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 18064 9976 18092 10016
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 20364 10053 20392 10084
rect 22066 10084 23704 10112
rect 20349 10047 20407 10053
rect 18196 10016 18241 10044
rect 19628 10016 20300 10044
rect 18196 10004 18202 10016
rect 19628 9976 19656 10016
rect 18064 9948 19656 9976
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9945 19763 9979
rect 20272 9976 20300 10016
rect 20349 10013 20361 10047
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 22066 9976 22094 10084
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 23014 10044 23020 10056
rect 22603 10016 23020 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 23676 10053 23704 10084
rect 24688 10084 25596 10112
rect 24578 10053 24584 10056
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 23891 10016 24409 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24545 10047 24584 10053
rect 24545 10013 24557 10047
rect 24545 10007 24584 10013
rect 20272 9948 22094 9976
rect 19705 9939 19763 9945
rect 16448 9880 17540 9908
rect 16448 9868 16454 9880
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18414 9908 18420 9920
rect 18104 9880 18420 9908
rect 18104 9868 18110 9880
rect 18414 9868 18420 9880
rect 18472 9908 18478 9920
rect 19720 9908 19748 9939
rect 22646 9936 22652 9988
rect 22704 9976 22710 9988
rect 22741 9979 22799 9985
rect 22741 9976 22753 9979
rect 22704 9948 22753 9976
rect 22704 9936 22710 9948
rect 22741 9945 22753 9948
rect 22787 9945 22799 9979
rect 22741 9939 22799 9945
rect 23584 9976 23612 10007
rect 23750 9976 23756 9988
rect 23584 9948 23756 9976
rect 18472 9880 19748 9908
rect 19797 9911 19855 9917
rect 18472 9868 18478 9880
rect 19797 9877 19809 9911
rect 19843 9908 19855 9911
rect 23584 9908 23612 9948
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 19843 9880 23612 9908
rect 24412 9908 24440 10007
rect 24578 10004 24584 10007
rect 24636 10004 24642 10056
rect 24688 10053 24716 10084
rect 25590 10072 25596 10084
rect 25648 10072 25654 10124
rect 25884 10112 25912 10143
rect 28442 10140 28448 10152
rect 28500 10140 28506 10192
rect 30929 10183 30987 10189
rect 30929 10149 30941 10183
rect 30975 10180 30987 10183
rect 31202 10180 31208 10192
rect 30975 10152 31208 10180
rect 30975 10149 30987 10152
rect 30929 10143 30987 10149
rect 31202 10140 31208 10152
rect 31260 10140 31266 10192
rect 26602 10112 26608 10124
rect 25700 10084 25912 10112
rect 26563 10084 26608 10112
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 24854 10004 24860 10056
rect 24912 10053 24918 10056
rect 24912 10047 24961 10053
rect 24912 10013 24915 10047
rect 24949 10013 24961 10047
rect 24912 10007 24961 10013
rect 24912 10004 24918 10007
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 25700 10044 25728 10084
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 30834 10112 30840 10124
rect 28368 10084 30840 10112
rect 25372 10016 25728 10044
rect 25777 10047 25835 10053
rect 25372 10004 25378 10016
rect 25777 10013 25789 10047
rect 25823 10013 25835 10047
rect 25777 10007 25835 10013
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9976 24823 9979
rect 25406 9976 25412 9988
rect 24811 9948 25412 9976
rect 24811 9945 24823 9948
rect 24765 9939 24823 9945
rect 25406 9936 25412 9948
rect 25464 9936 25470 9988
rect 24946 9908 24952 9920
rect 24412 9880 24952 9908
rect 19843 9877 19855 9880
rect 19797 9871 19855 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 25792 9908 25820 10007
rect 25866 10004 25872 10056
rect 25924 10044 25930 10056
rect 25961 10047 26019 10053
rect 25961 10044 25973 10047
rect 25924 10016 25973 10044
rect 25924 10004 25930 10016
rect 25961 10013 25973 10016
rect 26007 10013 26019 10047
rect 25961 10007 26019 10013
rect 26872 10047 26930 10053
rect 26872 10013 26884 10047
rect 26918 10044 26930 10047
rect 28368 10044 28396 10084
rect 30834 10072 30840 10084
rect 30892 10072 30898 10124
rect 31389 10115 31447 10121
rect 31389 10081 31401 10115
rect 31435 10112 31447 10115
rect 32490 10112 32496 10124
rect 31435 10084 32496 10112
rect 31435 10081 31447 10084
rect 31389 10075 31447 10081
rect 32490 10072 32496 10084
rect 32548 10072 32554 10124
rect 32950 10072 32956 10124
rect 33008 10112 33014 10124
rect 33502 10112 33508 10124
rect 33008 10084 33364 10112
rect 33463 10084 33508 10112
rect 33008 10072 33014 10084
rect 26918 10016 28396 10044
rect 26918 10013 26930 10016
rect 26872 10007 26930 10013
rect 28442 10004 28448 10056
rect 28500 10044 28506 10056
rect 28626 10044 28632 10056
rect 28500 10016 28545 10044
rect 28587 10016 28632 10044
rect 28500 10004 28506 10016
rect 28626 10004 28632 10016
rect 28684 10004 28690 10056
rect 29822 10004 29828 10056
rect 29880 10044 29886 10056
rect 30193 10047 30251 10053
rect 30193 10044 30205 10047
rect 29880 10016 30205 10044
rect 29880 10004 29886 10016
rect 30193 10013 30205 10016
rect 30239 10013 30251 10047
rect 30742 10044 30748 10056
rect 30703 10016 30748 10044
rect 30193 10007 30251 10013
rect 30742 10004 30748 10016
rect 30800 10004 30806 10056
rect 31573 10047 31631 10053
rect 31573 10013 31585 10047
rect 31619 10013 31631 10047
rect 31573 10007 31631 10013
rect 31757 10047 31815 10053
rect 31757 10013 31769 10047
rect 31803 10044 31815 10047
rect 32122 10044 32128 10056
rect 31803 10016 32128 10044
rect 31803 10013 31815 10016
rect 31757 10007 31815 10013
rect 26252 9948 28672 9976
rect 26050 9908 26056 9920
rect 25096 9880 25141 9908
rect 25792 9880 26056 9908
rect 25096 9868 25102 9880
rect 26050 9868 26056 9880
rect 26108 9908 26114 9920
rect 26252 9908 26280 9948
rect 26108 9880 26280 9908
rect 27985 9911 28043 9917
rect 26108 9868 26114 9880
rect 27985 9877 27997 9911
rect 28031 9908 28043 9911
rect 28442 9908 28448 9920
rect 28031 9880 28448 9908
rect 28031 9877 28043 9880
rect 27985 9871 28043 9877
rect 28442 9868 28448 9880
rect 28500 9868 28506 9920
rect 28644 9908 28672 9948
rect 29638 9936 29644 9988
rect 29696 9976 29702 9988
rect 29917 9979 29975 9985
rect 29917 9976 29929 9979
rect 29696 9948 29929 9976
rect 29696 9936 29702 9948
rect 29917 9945 29929 9948
rect 29963 9945 29975 9979
rect 31588 9976 31616 10007
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 32398 10044 32404 10056
rect 32359 10016 32404 10044
rect 32398 10004 32404 10016
rect 32456 10004 32462 10056
rect 33042 10044 33048 10056
rect 33003 10016 33048 10044
rect 33042 10004 33048 10016
rect 33100 10004 33106 10056
rect 33137 10047 33195 10053
rect 33137 10013 33149 10047
rect 33183 10044 33195 10047
rect 33226 10044 33232 10056
rect 33183 10016 33232 10044
rect 33183 10013 33195 10016
rect 33137 10007 33195 10013
rect 33226 10004 33232 10016
rect 33284 10004 33290 10056
rect 33336 10044 33364 10084
rect 33502 10072 33508 10084
rect 33560 10072 33566 10124
rect 33965 10047 34023 10053
rect 33965 10044 33977 10047
rect 33336 10016 33977 10044
rect 33965 10013 33977 10016
rect 34011 10013 34023 10047
rect 34146 10044 34152 10056
rect 34107 10016 34152 10044
rect 33965 10007 34023 10013
rect 34146 10004 34152 10016
rect 34204 10004 34210 10056
rect 34422 10004 34428 10056
rect 34480 10044 34486 10056
rect 35161 10047 35219 10053
rect 35161 10044 35173 10047
rect 34480 10016 35173 10044
rect 34480 10004 34486 10016
rect 35161 10013 35173 10016
rect 35207 10013 35219 10047
rect 35161 10007 35219 10013
rect 35897 10047 35955 10053
rect 35897 10013 35909 10047
rect 35943 10044 35955 10047
rect 36262 10044 36268 10056
rect 35943 10016 36268 10044
rect 35943 10013 35955 10016
rect 35897 10007 35955 10013
rect 29917 9939 29975 9945
rect 30024 9948 31616 9976
rect 30024 9908 30052 9948
rect 32030 9936 32036 9988
rect 32088 9976 32094 9988
rect 32861 9979 32919 9985
rect 32861 9976 32873 9979
rect 32088 9948 32873 9976
rect 32088 9936 32094 9948
rect 32861 9945 32873 9948
rect 32907 9945 32919 9979
rect 33778 9976 33784 9988
rect 32861 9939 32919 9945
rect 33336 9948 33784 9976
rect 28644 9880 30052 9908
rect 30101 9911 30159 9917
rect 30101 9877 30113 9911
rect 30147 9908 30159 9911
rect 30650 9908 30656 9920
rect 30147 9880 30656 9908
rect 30147 9877 30159 9880
rect 30101 9871 30159 9877
rect 30650 9868 30656 9880
rect 30708 9908 30714 9920
rect 31018 9908 31024 9920
rect 30708 9880 31024 9908
rect 30708 9868 30714 9880
rect 31018 9868 31024 9880
rect 31076 9868 31082 9920
rect 32214 9908 32220 9920
rect 32175 9880 32220 9908
rect 32214 9868 32220 9880
rect 32272 9868 32278 9920
rect 33134 9868 33140 9920
rect 33192 9908 33198 9920
rect 33336 9917 33364 9948
rect 33778 9936 33784 9948
rect 33836 9976 33842 9988
rect 35912 9976 35940 10007
rect 36262 10004 36268 10016
rect 36320 10004 36326 10056
rect 33836 9948 35940 9976
rect 33836 9936 33842 9948
rect 33321 9911 33379 9917
rect 33321 9908 33333 9911
rect 33192 9880 33333 9908
rect 33192 9868 33198 9880
rect 33321 9877 33333 9880
rect 33367 9877 33379 9911
rect 33321 9871 33379 9877
rect 33413 9911 33471 9917
rect 33413 9877 33425 9911
rect 33459 9908 33471 9911
rect 33594 9908 33600 9920
rect 33459 9880 33600 9908
rect 33459 9877 33471 9880
rect 33413 9871 33471 9877
rect 33594 9868 33600 9880
rect 33652 9868 33658 9920
rect 34054 9908 34060 9920
rect 34015 9880 34060 9908
rect 34054 9868 34060 9880
rect 34112 9868 34118 9920
rect 35253 9911 35311 9917
rect 35253 9877 35265 9911
rect 35299 9908 35311 9911
rect 35618 9908 35624 9920
rect 35299 9880 35624 9908
rect 35299 9877 35311 9880
rect 35253 9871 35311 9877
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 11330 9704 11336 9716
rect 2280 9676 11336 9704
rect 2280 9664 2286 9676
rect 11330 9664 11336 9676
rect 11388 9664 11394 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 16390 9704 16396 9716
rect 11664 9676 16396 9704
rect 11664 9664 11670 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 16724 9676 17233 9704
rect 16724 9664 16730 9676
rect 17221 9673 17233 9676
rect 17267 9673 17279 9707
rect 17221 9667 17279 9673
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21818 9704 21824 9716
rect 20772 9676 21824 9704
rect 20772 9664 20778 9676
rect 21818 9664 21824 9676
rect 21876 9704 21882 9716
rect 21876 9676 22784 9704
rect 21876 9664 21882 9676
rect 22756 9648 22784 9676
rect 23750 9664 23756 9716
rect 23808 9704 23814 9716
rect 24670 9704 24676 9716
rect 23808 9676 24676 9704
rect 23808 9664 23814 9676
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 25406 9704 25412 9716
rect 25367 9676 25412 9704
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 25590 9664 25596 9716
rect 25648 9704 25654 9716
rect 25648 9676 26280 9704
rect 25648 9664 25654 9676
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 4062 9636 4068 9648
rect 2188 9608 4068 9636
rect 2188 9596 2194 9608
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 4890 9636 4896 9648
rect 4448 9608 4896 9636
rect 4448 9577 4476 9608
rect 4890 9596 4896 9608
rect 4948 9636 4954 9648
rect 7006 9636 7012 9648
rect 4948 9608 7012 9636
rect 4948 9596 4954 9608
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 15657 9639 15715 9645
rect 7944 9608 12434 9636
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4700 9571 4758 9577
rect 4700 9537 4712 9571
rect 4746 9568 4758 9571
rect 5626 9568 5632 9580
rect 4746 9540 5632 9568
rect 4746 9537 4758 9540
rect 4700 9531 4758 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5776 9540 6377 9568
rect 5776 9528 5782 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6546 9568 6552 9580
rect 6507 9540 6552 9568
rect 6365 9531 6423 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6730 9568 6736 9580
rect 6687 9540 6736 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7834 9568 7840 9580
rect 7795 9540 7840 9568
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 6825 9435 6883 9441
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7944 9432 7972 9608
rect 8680 9577 8708 9608
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 8036 9500 8064 9531
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9364 9540 9781 9568
rect 9364 9528 9370 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10468 9540 10793 9568
rect 10468 9528 10474 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 11606 9568 11612 9580
rect 11567 9540 11612 9568
rect 10781 9531 10839 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 12406 9568 12434 9608
rect 15657 9605 15669 9639
rect 15703 9636 15715 9639
rect 16574 9636 16580 9648
rect 15703 9608 16580 9636
rect 15703 9605 15715 9608
rect 15657 9599 15715 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 18046 9636 18052 9648
rect 16776 9608 18052 9636
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12406 9540 13001 9568
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 8386 9500 8392 9512
rect 8036 9472 8392 9500
rect 8386 9460 8392 9472
rect 8444 9500 8450 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 8444 9472 8769 9500
rect 8444 9460 8450 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9500 9551 9503
rect 9674 9500 9680 9512
rect 9539 9472 9680 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 11790 9460 11796 9512
rect 11848 9500 11854 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11848 9472 11897 9500
rect 11848 9460 11854 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 13372 9500 13400 9531
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13596 9540 13737 9568
rect 13596 9528 13602 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14458 9568 14464 9580
rect 14415 9540 14464 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 11885 9463 11943 9469
rect 12406 9472 13400 9500
rect 6871 9404 7972 9432
rect 8205 9435 8263 9441
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 12406 9432 12434 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15344 9472 15761 9500
rect 15344 9460 15350 9472
rect 15749 9469 15761 9472
rect 15795 9500 15807 9503
rect 15838 9500 15844 9512
rect 15795 9472 15844 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 15948 9500 15976 9531
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16540 9540 16681 9568
rect 16540 9528 16546 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16776 9500 16804 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 18230 9645 18236 9648
rect 18224 9636 18236 9645
rect 18191 9608 18236 9636
rect 18224 9599 18236 9608
rect 18230 9596 18236 9599
rect 18288 9596 18294 9648
rect 22094 9636 22100 9648
rect 20456 9608 22100 9636
rect 20456 9580 20484 9608
rect 22094 9596 22100 9608
rect 22152 9596 22158 9648
rect 22738 9596 22744 9648
rect 22796 9596 22802 9648
rect 24302 9645 24308 9648
rect 24296 9636 24308 9645
rect 24263 9608 24308 9636
rect 24296 9599 24308 9608
rect 24302 9596 24308 9599
rect 24360 9596 24366 9648
rect 26252 9645 26280 9676
rect 29454 9664 29460 9716
rect 29512 9704 29518 9716
rect 31662 9704 31668 9716
rect 29512 9676 31668 9704
rect 29512 9664 29518 9676
rect 31662 9664 31668 9676
rect 31720 9664 31726 9716
rect 33502 9664 33508 9716
rect 33560 9704 33566 9716
rect 34517 9707 34575 9713
rect 34517 9704 34529 9707
rect 33560 9676 34529 9704
rect 33560 9664 33566 9676
rect 34517 9673 34529 9676
rect 34563 9704 34575 9707
rect 34563 9676 34744 9704
rect 34563 9673 34575 9676
rect 34517 9667 34575 9673
rect 26237 9639 26295 9645
rect 24504 9608 26096 9636
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 15948 9472 16804 9500
rect 16868 9500 16896 9531
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17083 9571 17141 9577
rect 17000 9540 17045 9568
rect 17000 9528 17006 9540
rect 17083 9537 17095 9571
rect 17129 9568 17141 9571
rect 17310 9568 17316 9580
rect 17129 9540 17316 9568
rect 17129 9537 17141 9540
rect 17083 9531 17141 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 20349 9571 20407 9577
rect 17788 9540 19334 9568
rect 17218 9500 17224 9512
rect 16868 9472 17224 9500
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 8251 9404 12434 9432
rect 13173 9435 13231 9441
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 17788 9432 17816 9540
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 17957 9503 18015 9509
rect 17957 9500 17969 9503
rect 17920 9472 17969 9500
rect 17920 9460 17926 9472
rect 17957 9469 17969 9472
rect 18003 9469 18015 9503
rect 19306 9500 19334 9540
rect 20349 9537 20361 9571
rect 20395 9568 20407 9571
rect 20438 9568 20444 9580
rect 20395 9540 20444 9568
rect 20395 9537 20407 9540
rect 20349 9531 20407 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 20714 9568 20720 9580
rect 20579 9540 20720 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 20548 9500 20576 9531
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 20990 9568 20996 9580
rect 20951 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9568 22247 9571
rect 22278 9568 22284 9580
rect 22235 9540 22284 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 22462 9577 22468 9580
rect 22456 9531 22468 9577
rect 22520 9568 22526 9580
rect 24026 9568 24032 9580
rect 22520 9540 22556 9568
rect 23987 9540 24032 9568
rect 22462 9528 22468 9531
rect 22520 9528 22526 9540
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24504 9568 24532 9608
rect 26068 9580 26096 9608
rect 26237 9605 26249 9639
rect 26283 9636 26295 9639
rect 26786 9636 26792 9648
rect 26283 9608 26792 9636
rect 26283 9605 26295 9608
rect 26237 9599 26295 9605
rect 26786 9596 26792 9608
rect 26844 9596 26850 9648
rect 29086 9596 29092 9648
rect 29144 9636 29150 9648
rect 30009 9639 30067 9645
rect 30009 9636 30021 9639
rect 29144 9608 30021 9636
rect 29144 9596 29150 9608
rect 30009 9605 30021 9608
rect 30055 9605 30067 9639
rect 30009 9599 30067 9605
rect 30116 9608 31754 9636
rect 24136 9540 24532 9568
rect 19306 9472 20576 9500
rect 17957 9463 18015 9469
rect 23750 9460 23756 9512
rect 23808 9500 23814 9512
rect 24136 9500 24164 9540
rect 24854 9528 24860 9580
rect 24912 9568 24918 9580
rect 25866 9568 25872 9580
rect 24912 9540 25872 9568
rect 24912 9528 24918 9540
rect 25866 9528 25872 9540
rect 25924 9528 25930 9580
rect 26050 9568 26056 9580
rect 26011 9540 26056 9568
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 26973 9571 27031 9577
rect 26973 9568 26985 9571
rect 26160 9540 26985 9568
rect 23808 9472 24164 9500
rect 23808 9460 23814 9472
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 26160 9500 26188 9540
rect 26973 9537 26985 9540
rect 27019 9537 27031 9571
rect 27154 9568 27160 9580
rect 27115 9540 27160 9568
rect 26973 9531 27031 9537
rect 27154 9528 27160 9540
rect 27212 9528 27218 9580
rect 27976 9571 28034 9577
rect 27976 9537 27988 9571
rect 28022 9568 28034 9571
rect 30116 9568 30144 9608
rect 28022 9540 30144 9568
rect 30193 9571 30251 9577
rect 28022 9537 28034 9540
rect 27976 9531 28034 9537
rect 30193 9537 30205 9571
rect 30239 9568 30251 9571
rect 30745 9571 30803 9577
rect 30745 9568 30757 9571
rect 30239 9540 30757 9568
rect 30239 9537 30251 9540
rect 30193 9531 30251 9537
rect 30745 9537 30757 9540
rect 30791 9568 30803 9571
rect 31018 9568 31024 9580
rect 30791 9540 31024 9568
rect 30791 9537 30803 9540
rect 30745 9531 30803 9537
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9537 31447 9571
rect 31570 9568 31576 9580
rect 31531 9540 31576 9568
rect 31389 9531 31447 9537
rect 25280 9472 26188 9500
rect 25280 9460 25286 9472
rect 26602 9460 26608 9512
rect 26660 9500 26666 9512
rect 27709 9503 27767 9509
rect 27709 9500 27721 9503
rect 26660 9472 27721 9500
rect 26660 9460 26666 9472
rect 27709 9469 27721 9472
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 19702 9432 19708 9444
rect 13219 9404 17816 9432
rect 19260 9404 19708 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5859 9336 6377 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 6365 9333 6377 9336
rect 6411 9364 6423 9367
rect 6454 9364 6460 9376
rect 6411 9336 6460 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 7984 9336 8677 9364
rect 7984 9324 7990 9336
rect 8665 9333 8677 9336
rect 8711 9333 8723 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 8665 9327 8723 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10873 9367 10931 9373
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 11974 9364 11980 9376
rect 10919 9336 11980 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 15378 9364 15384 9376
rect 12216 9336 15384 9364
rect 12216 9324 12222 9336
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 19260 9364 19288 9404
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20622 9432 20628 9444
rect 20036 9404 20628 9432
rect 20036 9392 20042 9404
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 21082 9432 21088 9444
rect 21043 9404 21088 9432
rect 21082 9392 21088 9404
rect 21140 9392 21146 9444
rect 28718 9392 28724 9444
rect 28776 9432 28782 9444
rect 31404 9432 31432 9531
rect 31570 9528 31576 9540
rect 31628 9528 31634 9580
rect 31726 9568 31754 9608
rect 32214 9596 32220 9648
rect 32272 9636 32278 9648
rect 32370 9639 32428 9645
rect 32370 9636 32382 9639
rect 32272 9608 32382 9636
rect 32272 9596 32278 9608
rect 32370 9605 32382 9608
rect 32416 9605 32428 9639
rect 34606 9636 34612 9648
rect 32370 9599 32428 9605
rect 32508 9608 34612 9636
rect 32508 9568 32536 9608
rect 34606 9596 34612 9608
rect 34664 9596 34670 9648
rect 34716 9636 34744 9676
rect 34716 9608 35296 9636
rect 34238 9568 34244 9580
rect 31726 9540 32536 9568
rect 34199 9540 34244 9568
rect 34238 9528 34244 9540
rect 34296 9528 34302 9580
rect 35268 9577 35296 9608
rect 34379 9571 34437 9577
rect 34379 9537 34391 9571
rect 34425 9568 34437 9571
rect 35069 9571 35127 9577
rect 35069 9568 35081 9571
rect 34425 9540 34560 9568
rect 34425 9537 34437 9540
rect 34379 9531 34437 9537
rect 31846 9460 31852 9512
rect 31904 9500 31910 9512
rect 32125 9503 32183 9509
rect 32125 9500 32137 9503
rect 31904 9472 32137 9500
rect 31904 9460 31910 9472
rect 32125 9469 32137 9472
rect 32171 9469 32183 9503
rect 32125 9463 32183 9469
rect 33870 9460 33876 9512
rect 33928 9500 33934 9512
rect 34149 9503 34207 9509
rect 34149 9500 34161 9503
rect 33928 9472 34161 9500
rect 33928 9460 33934 9472
rect 34149 9469 34161 9472
rect 34195 9469 34207 9503
rect 34149 9463 34207 9469
rect 28776 9404 31432 9432
rect 34532 9432 34560 9540
rect 34624 9540 35081 9568
rect 34624 9512 34652 9540
rect 35069 9537 35081 9540
rect 35115 9537 35127 9571
rect 35069 9531 35127 9537
rect 35253 9571 35311 9577
rect 35253 9537 35265 9571
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 35345 9571 35403 9577
rect 35345 9537 35357 9571
rect 35391 9568 35403 9571
rect 35618 9568 35624 9580
rect 35391 9540 35624 9568
rect 35391 9537 35403 9540
rect 35345 9531 35403 9537
rect 35618 9528 35624 9540
rect 35676 9528 35682 9580
rect 35805 9571 35863 9577
rect 35805 9537 35817 9571
rect 35851 9537 35863 9571
rect 35986 9568 35992 9580
rect 35947 9540 35992 9568
rect 35805 9531 35863 9537
rect 34606 9460 34612 9512
rect 34664 9500 34670 9512
rect 34664 9472 34709 9500
rect 34664 9460 34670 9472
rect 35434 9460 35440 9512
rect 35492 9500 35498 9512
rect 35820 9500 35848 9531
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 35492 9472 35848 9500
rect 35492 9460 35498 9472
rect 34790 9432 34796 9444
rect 34532 9404 34796 9432
rect 28776 9392 28782 9404
rect 34790 9392 34796 9404
rect 34848 9392 34854 9444
rect 16163 9336 19288 9364
rect 19337 9367 19395 9373
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19426 9364 19432 9376
rect 19383 9336 19432 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 21910 9324 21916 9376
rect 21968 9364 21974 9376
rect 23569 9367 23627 9373
rect 23569 9364 23581 9367
rect 21968 9336 23581 9364
rect 21968 9324 21974 9336
rect 23569 9333 23581 9336
rect 23615 9333 23627 9367
rect 23569 9327 23627 9333
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 26973 9367 27031 9373
rect 26973 9364 26985 9367
rect 25464 9336 26985 9364
rect 25464 9324 25470 9336
rect 26973 9333 26985 9336
rect 27019 9333 27031 9367
rect 26973 9327 27031 9333
rect 29089 9367 29147 9373
rect 29089 9333 29101 9367
rect 29135 9364 29147 9367
rect 29178 9364 29184 9376
rect 29135 9336 29184 9364
rect 29135 9333 29147 9336
rect 29089 9327 29147 9333
rect 29178 9324 29184 9336
rect 29236 9324 29242 9376
rect 29638 9324 29644 9376
rect 29696 9364 29702 9376
rect 30837 9367 30895 9373
rect 30837 9364 30849 9367
rect 29696 9336 30849 9364
rect 29696 9324 29702 9336
rect 30837 9333 30849 9336
rect 30883 9333 30895 9367
rect 30837 9327 30895 9333
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 31389 9367 31447 9373
rect 31389 9364 31401 9367
rect 31168 9336 31401 9364
rect 31168 9324 31174 9336
rect 31389 9333 31401 9336
rect 31435 9333 31447 9367
rect 31389 9327 31447 9333
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 33042 9364 33048 9376
rect 31812 9336 33048 9364
rect 31812 9324 31818 9336
rect 33042 9324 33048 9336
rect 33100 9364 33106 9376
rect 33505 9367 33563 9373
rect 33505 9364 33517 9367
rect 33100 9336 33517 9364
rect 33100 9324 33106 9336
rect 33505 9333 33517 9336
rect 33551 9364 33563 9367
rect 33870 9364 33876 9376
rect 33551 9336 33876 9364
rect 33551 9333 33563 9336
rect 33505 9327 33563 9333
rect 33870 9324 33876 9336
rect 33928 9324 33934 9376
rect 33965 9367 34023 9373
rect 33965 9333 33977 9367
rect 34011 9364 34023 9367
rect 34146 9364 34152 9376
rect 34011 9336 34152 9364
rect 34011 9333 34023 9336
rect 33965 9327 34023 9333
rect 34146 9324 34152 9336
rect 34204 9324 34210 9376
rect 34514 9324 34520 9376
rect 34572 9364 34578 9376
rect 35161 9367 35219 9373
rect 35161 9364 35173 9367
rect 34572 9336 35173 9364
rect 34572 9324 34578 9336
rect 35161 9333 35173 9336
rect 35207 9333 35219 9367
rect 35802 9364 35808 9376
rect 35763 9336 35808 9364
rect 35161 9327 35219 9333
rect 35802 9324 35808 9336
rect 35860 9324 35866 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5718 9160 5724 9172
rect 4120 9132 5580 9160
rect 5679 9132 5724 9160
rect 4120 9120 4126 9132
rect 5552 9092 5580 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 8018 9160 8024 9172
rect 7979 9132 8024 9160
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8386 9160 8392 9172
rect 8347 9132 8392 9160
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 10410 9160 10416 9172
rect 8956 9132 10416 9160
rect 8956 9092 8984 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10594 9160 10600 9172
rect 10555 9132 10600 9160
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12066 9160 12072 9172
rect 12023 9132 12072 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 13538 9160 13544 9172
rect 13499 9132 13544 9160
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9129 14151 9163
rect 14093 9123 14151 9129
rect 14461 9163 14519 9169
rect 14461 9129 14473 9163
rect 14507 9160 14519 9163
rect 15286 9160 15292 9172
rect 14507 9132 15292 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 5552 9064 8984 9092
rect 9030 9052 9036 9104
rect 9088 9092 9094 9104
rect 14108 9092 14136 9123
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 16025 9163 16083 9169
rect 16025 9160 16037 9163
rect 15436 9132 16037 9160
rect 15436 9120 15442 9132
rect 16025 9129 16037 9132
rect 16071 9129 16083 9163
rect 18874 9160 18880 9172
rect 16025 9123 16083 9129
rect 16684 9132 18880 9160
rect 9088 9064 11928 9092
rect 9088 9052 9094 9064
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6638 8984 6644 8996
rect 6696 9024 6702 9036
rect 6696 8996 7696 9024
rect 6696 8984 6702 8996
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4890 8956 4896 8968
rect 4387 8928 4896 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6328 8928 6377 8956
rect 6328 8916 6334 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6733 8959 6791 8965
rect 6512 8928 6557 8956
rect 6512 8916 6518 8928
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7466 8956 7472 8968
rect 7423 8928 7472 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 4614 8897 4620 8900
rect 4608 8851 4620 8897
rect 4672 8888 4678 8900
rect 4672 8860 4708 8888
rect 4614 8848 4620 8851
rect 4672 8848 4678 8860
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 6748 8888 6776 8919
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7668 8956 7696 8996
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7800 8996 8033 9024
rect 7800 8984 7806 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8812 8996 9505 9024
rect 8812 8984 8818 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 11054 9024 11060 9036
rect 9493 8987 9551 8993
rect 9600 8996 11060 9024
rect 8205 8959 8263 8965
rect 7668 8928 8156 8956
rect 5500 8860 6776 8888
rect 5500 8848 5506 8860
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 7929 8891 7987 8897
rect 7929 8888 7941 8891
rect 6880 8860 7941 8888
rect 6880 8848 6886 8860
rect 7929 8857 7941 8860
rect 7975 8857 7987 8891
rect 8128 8888 8156 8928
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8570 8956 8576 8968
rect 8251 8928 8576 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8570 8916 8576 8928
rect 8628 8956 8634 8968
rect 8938 8956 8944 8968
rect 8628 8928 8944 8956
rect 8628 8916 8634 8928
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9600 8888 9628 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11388 8996 11836 9024
rect 11388 8984 11394 8996
rect 11808 8968 11836 8996
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11238 8956 11244 8968
rect 11195 8928 11244 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 8128 8860 9628 8888
rect 7929 8851 7987 8857
rect 7190 8820 7196 8832
rect 7151 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10796 8820 10824 8919
rect 10888 8888 10916 8919
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11572 8928 11621 8956
rect 11572 8916 11578 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 11609 8919 11667 8925
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 11422 8888 11428 8900
rect 10888 8860 11428 8888
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11900 8888 11928 9064
rect 13188 9064 14136 9092
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 12032 8928 12449 8956
rect 12032 8916 12038 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 11900 8860 12756 8888
rect 10962 8820 10968 8832
rect 9824 8792 10968 8820
rect 9824 8780 9830 8792
rect 10962 8780 10968 8792
rect 11020 8820 11026 8832
rect 12066 8820 12072 8832
rect 11020 8792 12072 8820
rect 11020 8780 11026 8792
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12526 8820 12532 8832
rect 12400 8792 12532 8820
rect 12400 8780 12406 8792
rect 12526 8780 12532 8792
rect 12584 8820 12590 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12584 8792 12633 8820
rect 12584 8780 12590 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 12728 8820 12756 8860
rect 12894 8848 12900 8900
rect 12952 8888 12958 8900
rect 13188 8897 13216 9064
rect 15746 9052 15752 9104
rect 15804 9092 15810 9104
rect 16684 9092 16712 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 19889 9163 19947 9169
rect 19889 9129 19901 9163
rect 19935 9160 19947 9163
rect 20162 9160 20168 9172
rect 19935 9132 20168 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 20162 9120 20168 9132
rect 20220 9160 20226 9172
rect 20806 9160 20812 9172
rect 20220 9132 20812 9160
rect 20220 9120 20226 9132
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 22066 9132 23520 9160
rect 15804 9064 16712 9092
rect 15804 9052 15810 9064
rect 18322 9052 18328 9104
rect 18380 9092 18386 9104
rect 20990 9092 20996 9104
rect 18380 9064 20996 9092
rect 18380 9052 18386 9064
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 15177 9027 15235 9033
rect 13412 8996 14136 9024
rect 13412 8984 13418 8996
rect 13372 8956 13400 8984
rect 14108 8965 14136 8996
rect 15177 8993 15189 9027
rect 15223 9024 15235 9027
rect 19610 9024 19616 9036
rect 15223 8996 16068 9024
rect 15223 8993 15235 8996
rect 15177 8987 15235 8993
rect 13280 8928 13400 8956
rect 14093 8959 14151 8965
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12952 8860 13185 8888
rect 12952 8848 12958 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 13280 8820 13308 8928
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 14093 8919 14151 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15378 8956 15384 8968
rect 15339 8928 15384 8956
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15896 8928 15945 8956
rect 15896 8916 15902 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 14292 8888 14320 8916
rect 13403 8860 14320 8888
rect 15105 8891 15163 8897
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 15105 8857 15117 8891
rect 15151 8888 15163 8891
rect 16040 8888 16068 8996
rect 18524 8996 19616 9024
rect 16669 8959 16727 8965
rect 16669 8925 16681 8959
rect 16715 8956 16727 8959
rect 16758 8956 16764 8968
rect 16715 8928 16764 8956
rect 16715 8925 16727 8928
rect 16669 8919 16727 8925
rect 16758 8916 16764 8928
rect 16816 8956 16822 8968
rect 17862 8956 17868 8968
rect 16816 8928 17868 8956
rect 16816 8916 16822 8928
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18524 8965 18552 8996
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 19150 8956 19156 8968
rect 18739 8928 19156 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19260 8965 19288 8996
rect 19610 8984 19616 8996
rect 19668 8984 19674 9036
rect 20364 9024 20392 9064
rect 20990 9052 20996 9064
rect 21048 9092 21054 9104
rect 22066 9092 22094 9132
rect 21048 9064 22094 9092
rect 23492 9092 23520 9132
rect 23566 9120 23572 9172
rect 23624 9160 23630 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23624 9132 23673 9160
rect 23624 9120 23630 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 26326 9160 26332 9172
rect 24820 9132 26332 9160
rect 24820 9120 24826 9132
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 28810 9120 28816 9172
rect 28868 9160 28874 9172
rect 31754 9160 31760 9172
rect 28868 9132 31760 9160
rect 28868 9120 28874 9132
rect 31754 9120 31760 9132
rect 31812 9120 31818 9172
rect 32030 9160 32036 9172
rect 31991 9132 32036 9160
rect 32030 9120 32036 9132
rect 32088 9120 32094 9172
rect 32217 9163 32275 9169
rect 32217 9129 32229 9163
rect 32263 9160 32275 9163
rect 32398 9160 32404 9172
rect 32263 9132 32404 9160
rect 32263 9129 32275 9132
rect 32217 9123 32275 9129
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 33594 9120 33600 9172
rect 33652 9160 33658 9172
rect 33965 9163 34023 9169
rect 33965 9160 33977 9163
rect 33652 9132 33977 9160
rect 33652 9120 33658 9132
rect 33965 9129 33977 9132
rect 34011 9129 34023 9163
rect 33965 9123 34023 9129
rect 34149 9163 34207 9169
rect 34149 9129 34161 9163
rect 34195 9160 34207 9163
rect 34606 9160 34612 9172
rect 34195 9132 34612 9160
rect 34195 9129 34207 9132
rect 34149 9123 34207 9129
rect 34606 9120 34612 9132
rect 34664 9120 34670 9172
rect 35802 9160 35808 9172
rect 34716 9132 35808 9160
rect 24854 9092 24860 9104
rect 23492 9064 24860 9092
rect 21048 9052 21054 9064
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 26344 9092 26372 9120
rect 28166 9092 28172 9104
rect 26344 9064 28172 9092
rect 28166 9052 28172 9064
rect 28224 9052 28230 9104
rect 28718 9052 28724 9104
rect 28776 9092 28782 9104
rect 28776 9064 28821 9092
rect 28776 9052 28782 9064
rect 33042 9052 33048 9104
rect 33100 9092 33106 9104
rect 33318 9092 33324 9104
rect 33100 9064 33324 9092
rect 33100 9052 33106 9064
rect 33318 9052 33324 9064
rect 33376 9052 33382 9104
rect 33410 9052 33416 9104
rect 33468 9092 33474 9104
rect 34716 9092 34744 9132
rect 35802 9120 35808 9132
rect 35860 9120 35866 9172
rect 33468 9064 34744 9092
rect 33468 9052 33474 9064
rect 20272 8996 20392 9024
rect 19245 8959 19303 8965
rect 19245 8925 19257 8959
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 19978 8956 19984 8968
rect 19475 8928 19984 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20162 8965 20168 8968
rect 20119 8959 20168 8965
rect 20119 8925 20131 8959
rect 20165 8925 20168 8959
rect 20119 8919 20168 8925
rect 20162 8916 20168 8919
rect 20220 8916 20226 8968
rect 20272 8965 20300 8996
rect 21082 8984 21088 9036
rect 21140 9024 21146 9036
rect 22278 9024 22284 9036
rect 21140 8996 22094 9024
rect 22191 8996 22284 9024
rect 21140 8984 21146 8996
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20346 8916 20352 8968
rect 20404 8956 20410 8968
rect 21192 8965 21220 8996
rect 20533 8959 20591 8965
rect 20404 8928 20449 8956
rect 20404 8916 20410 8928
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 21177 8959 21235 8965
rect 21177 8956 21189 8959
rect 20579 8928 21189 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 21177 8925 21189 8928
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21324 8928 21373 8956
rect 21324 8916 21330 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 16914 8891 16972 8897
rect 16914 8888 16926 8891
rect 15151 8860 15976 8888
rect 16040 8860 16926 8888
rect 15151 8857 15163 8860
rect 15105 8851 15163 8857
rect 15286 8820 15292 8832
rect 12728 8792 13308 8820
rect 15247 8792 15292 8820
rect 12621 8783 12679 8789
rect 15286 8780 15292 8792
rect 15344 8820 15350 8832
rect 15746 8820 15752 8832
rect 15344 8792 15752 8820
rect 15344 8780 15350 8792
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 15948 8820 15976 8860
rect 16914 8857 16926 8860
rect 16960 8857 16972 8891
rect 16914 8851 16972 8857
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8857 18659 8891
rect 19886 8888 19892 8900
rect 18601 8851 18659 8857
rect 19260 8860 19892 8888
rect 17586 8820 17592 8832
rect 15948 8792 17592 8820
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18616 8820 18644 8851
rect 19260 8820 19288 8860
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 21468 8888 21496 8919
rect 20496 8860 21496 8888
rect 22066 8888 22094 8996
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 24026 8984 24032 9036
rect 24084 9024 24090 9036
rect 24949 9027 25007 9033
rect 24949 9024 24961 9027
rect 24084 8996 24961 9024
rect 24084 8984 24090 8996
rect 24949 8993 24961 8996
rect 24995 8993 25007 9027
rect 24949 8987 25007 8993
rect 26142 8984 26148 9036
rect 26200 8984 26206 9036
rect 26786 9024 26792 9036
rect 26747 8996 26792 9024
rect 26786 8984 26792 8996
rect 26844 8984 26850 9036
rect 28184 9024 28212 9052
rect 29638 9024 29644 9036
rect 28184 8996 28585 9024
rect 29599 8996 29644 9024
rect 22296 8956 22324 8984
rect 24044 8956 24072 8984
rect 22296 8928 24072 8956
rect 25216 8959 25274 8965
rect 25216 8925 25228 8959
rect 25262 8956 25274 8959
rect 26160 8956 26188 8984
rect 25262 8928 26188 8956
rect 25262 8925 25274 8928
rect 25216 8919 25274 8925
rect 26694 8916 26700 8968
rect 26752 8956 26758 8968
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 26752 8928 27077 8956
rect 26752 8916 26758 8928
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 22278 8888 22284 8900
rect 22066 8860 22284 8888
rect 20496 8848 20502 8860
rect 22278 8848 22284 8860
rect 22336 8848 22342 8900
rect 22554 8897 22560 8900
rect 22548 8888 22560 8897
rect 22515 8860 22560 8888
rect 22548 8851 22560 8860
rect 22554 8848 22560 8851
rect 22612 8848 22618 8900
rect 22738 8848 22744 8900
rect 22796 8888 22802 8900
rect 27080 8888 27108 8919
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 28258 8965 28264 8968
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 27580 8928 28089 8956
rect 27580 8916 27586 8928
rect 28077 8925 28089 8928
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 28225 8959 28264 8965
rect 28225 8925 28237 8959
rect 28225 8919 28264 8925
rect 28258 8916 28264 8919
rect 28316 8916 28322 8968
rect 28442 8956 28448 8968
rect 28403 8928 28448 8956
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 28557 8965 28585 8996
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 34054 9024 34060 9036
rect 31726 8996 34060 9024
rect 28542 8959 28600 8965
rect 28542 8925 28554 8959
rect 28588 8925 28600 8959
rect 28542 8919 28600 8925
rect 29908 8959 29966 8965
rect 29908 8925 29920 8959
rect 29954 8956 29966 8959
rect 31726 8956 31754 8996
rect 34054 8984 34060 8996
rect 34112 8984 34118 9036
rect 29954 8928 31754 8956
rect 29954 8925 29966 8928
rect 29908 8919 29966 8925
rect 32214 8916 32220 8968
rect 32272 8956 32278 8968
rect 32861 8959 32919 8965
rect 32861 8956 32873 8959
rect 32272 8928 32873 8956
rect 32272 8916 32278 8928
rect 32861 8925 32873 8928
rect 32907 8925 32919 8959
rect 32861 8919 32919 8925
rect 32953 8959 33011 8965
rect 32953 8925 32965 8959
rect 32999 8956 33011 8959
rect 33226 8956 33232 8968
rect 32999 8928 33232 8956
rect 32999 8925 33011 8928
rect 32953 8919 33011 8925
rect 33226 8916 33232 8928
rect 33284 8916 33290 8968
rect 33321 8959 33379 8965
rect 33321 8925 33333 8959
rect 33367 8956 33379 8959
rect 33502 8956 33508 8968
rect 33367 8928 33508 8956
rect 33367 8925 33379 8928
rect 33321 8919 33379 8925
rect 33502 8916 33508 8928
rect 33560 8916 33566 8968
rect 34514 8956 34520 8968
rect 33704 8928 34520 8956
rect 28353 8891 28411 8897
rect 28353 8888 28365 8891
rect 22796 8860 27016 8888
rect 27080 8860 28365 8888
rect 22796 8848 22802 8860
rect 18616 8792 19288 8820
rect 19337 8823 19395 8829
rect 19337 8789 19349 8823
rect 19383 8820 19395 8823
rect 19426 8820 19432 8832
rect 19383 8792 19432 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 20993 8823 21051 8829
rect 20993 8820 21005 8823
rect 20404 8792 21005 8820
rect 20404 8780 20410 8792
rect 20993 8789 21005 8792
rect 21039 8789 21051 8823
rect 20993 8783 21051 8789
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 25222 8820 25228 8832
rect 22428 8792 25228 8820
rect 22428 8780 22434 8792
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 25314 8780 25320 8832
rect 25372 8820 25378 8832
rect 25866 8820 25872 8832
rect 25372 8792 25872 8820
rect 25372 8780 25378 8792
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 26329 8823 26387 8829
rect 26329 8820 26341 8823
rect 26016 8792 26341 8820
rect 26016 8780 26022 8792
rect 26329 8789 26341 8792
rect 26375 8789 26387 8823
rect 26988 8820 27016 8860
rect 28353 8857 28365 8860
rect 28399 8888 28411 8891
rect 28902 8888 28908 8900
rect 28399 8860 28908 8888
rect 28399 8857 28411 8860
rect 28353 8851 28411 8857
rect 28902 8848 28908 8860
rect 28960 8848 28966 8900
rect 30742 8888 30748 8900
rect 30392 8860 30748 8888
rect 30392 8820 30420 8860
rect 30742 8848 30748 8860
rect 30800 8848 30806 8900
rect 31849 8891 31907 8897
rect 31849 8857 31861 8891
rect 31895 8888 31907 8891
rect 32306 8888 32312 8900
rect 31895 8860 32312 8888
rect 31895 8857 31907 8860
rect 31849 8851 31907 8857
rect 32306 8848 32312 8860
rect 32364 8848 32370 8900
rect 33704 8888 33732 8928
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 34698 8956 34704 8968
rect 34659 8928 34704 8956
rect 34698 8916 34704 8928
rect 34756 8916 34762 8968
rect 32508 8860 33732 8888
rect 26988 8792 30420 8820
rect 26329 8783 26387 8789
rect 30466 8780 30472 8832
rect 30524 8820 30530 8832
rect 31021 8823 31079 8829
rect 31021 8820 31033 8823
rect 30524 8792 31033 8820
rect 30524 8780 30530 8792
rect 31021 8789 31033 8792
rect 31067 8789 31079 8823
rect 31021 8783 31079 8789
rect 32059 8823 32117 8829
rect 32059 8789 32071 8823
rect 32105 8820 32117 8823
rect 32508 8820 32536 8860
rect 33778 8848 33784 8900
rect 33836 8888 33842 8900
rect 33836 8860 33881 8888
rect 33836 8848 33842 8860
rect 33962 8848 33968 8900
rect 34020 8897 34026 8900
rect 34020 8891 34039 8897
rect 34027 8857 34039 8891
rect 34020 8851 34039 8857
rect 34020 8848 34026 8851
rect 34422 8848 34428 8900
rect 34480 8888 34486 8900
rect 34946 8891 35004 8897
rect 34946 8888 34958 8891
rect 34480 8860 34958 8888
rect 34480 8848 34486 8860
rect 34946 8857 34958 8860
rect 34992 8857 35004 8891
rect 34946 8851 35004 8857
rect 32674 8820 32680 8832
rect 32105 8792 32536 8820
rect 32635 8792 32680 8820
rect 32105 8789 32117 8792
rect 32059 8783 32117 8789
rect 32674 8780 32680 8792
rect 32732 8780 32738 8832
rect 33134 8820 33140 8832
rect 33095 8792 33140 8820
rect 33134 8780 33140 8792
rect 33192 8780 33198 8832
rect 33229 8823 33287 8829
rect 33229 8789 33241 8823
rect 33275 8820 33287 8823
rect 33594 8820 33600 8832
rect 33275 8792 33600 8820
rect 33275 8789 33287 8792
rect 33229 8783 33287 8789
rect 33594 8780 33600 8792
rect 33652 8780 33658 8832
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 36081 8823 36139 8829
rect 36081 8820 36093 8823
rect 34848 8792 36093 8820
rect 34848 8780 34854 8792
rect 36081 8789 36093 8792
rect 36127 8789 36139 8823
rect 36081 8783 36139 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 4614 8616 4620 8628
rect 4575 8588 4620 8616
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5684 8588 6377 8616
rect 5684 8576 5690 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 8938 8616 8944 8628
rect 8899 8588 8944 8616
rect 6365 8579 6423 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 16298 8616 16304 8628
rect 9272 8588 16304 8616
rect 9272 8576 9278 8588
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 17000 8588 19932 8616
rect 17000 8576 17006 8588
rect 19904 8560 19932 8588
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20220 8588 21189 8616
rect 20220 8576 20226 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 24121 8619 24179 8625
rect 24121 8616 24133 8619
rect 21784 8588 24133 8616
rect 21784 8576 21790 8588
rect 24121 8585 24133 8588
rect 24167 8585 24179 8619
rect 27246 8616 27252 8628
rect 24121 8579 24179 8585
rect 25884 8588 27252 8616
rect 6270 8548 6276 8560
rect 5460 8520 6276 8548
rect 5460 8489 5488 8520
rect 6270 8508 6276 8520
rect 6328 8548 6334 8560
rect 6730 8548 6736 8560
rect 6328 8520 6736 8548
rect 6328 8508 6334 8520
rect 6730 8508 6736 8520
rect 6788 8548 6794 8560
rect 9766 8548 9772 8560
rect 6788 8520 9772 8548
rect 6788 8508 6794 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 10560 8520 12434 8548
rect 10560 8508 10566 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5718 8480 5724 8492
rect 5583 8452 5724 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 4816 8344 4844 8443
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5828 8412 5856 8443
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6420 8452 6561 8480
rect 6420 8440 6426 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7834 8489 7840 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7064 8452 7573 8480
rect 7064 8440 7070 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7828 8443 7840 8489
rect 7892 8480 7898 8492
rect 9398 8480 9404 8492
rect 7892 8452 7928 8480
rect 9359 8452 9404 8480
rect 7834 8440 7840 8443
rect 7892 8440 7898 8452
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9582 8480 9588 8492
rect 9543 8452 9588 8480
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 11885 8483 11943 8489
rect 10459 8452 11468 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 11330 8412 11336 8424
rect 5132 8384 5856 8412
rect 8588 8384 11336 8412
rect 5132 8372 5138 8384
rect 5534 8344 5540 8356
rect 4816 8316 5540 8344
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 6638 8344 6644 8356
rect 5767 8316 6644 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 8588 8344 8616 8384
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 8496 8316 8616 8344
rect 5258 8276 5264 8288
rect 5219 8248 5264 8276
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 7282 8276 7288 8288
rect 5408 8248 7288 8276
rect 5408 8236 5414 8248
rect 7282 8236 7288 8248
rect 7340 8276 7346 8288
rect 8496 8276 8524 8316
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9769 8347 9827 8353
rect 9769 8344 9781 8347
rect 8720 8316 9781 8344
rect 8720 8304 8726 8316
rect 9769 8313 9781 8316
rect 9815 8313 9827 8347
rect 11440 8344 11468 8452
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 11885 8443 11943 8449
rect 11900 8412 11928 8443
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12406 8480 12434 8520
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 14645 8551 14703 8557
rect 14645 8548 14657 8551
rect 13780 8520 14657 8548
rect 13780 8508 13786 8520
rect 14645 8517 14657 8520
rect 14691 8517 14703 8551
rect 14645 8511 14703 8517
rect 14743 8520 18828 8548
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12406 8452 12541 8480
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 13354 8480 13360 8492
rect 13315 8452 13360 8480
rect 12529 8443 12587 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 14458 8480 14464 8492
rect 14419 8452 14464 8480
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 13372 8412 13400 8440
rect 11900 8384 13400 8412
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 14743 8412 14771 8520
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15470 8480 15476 8492
rect 15335 8452 15476 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16482 8480 16488 8492
rect 15611 8452 16488 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17175 8452 17693 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17681 8449 17693 8452
rect 17727 8480 17739 8483
rect 17954 8480 17960 8492
rect 17727 8452 17960 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18800 8489 18828 8520
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 19490 8551 19548 8557
rect 19490 8548 19502 8551
rect 19392 8520 19502 8548
rect 19392 8508 19398 8520
rect 19490 8517 19502 8520
rect 19536 8517 19548 8551
rect 19490 8511 19548 8517
rect 19886 8508 19892 8560
rect 19944 8508 19950 8560
rect 22005 8551 22063 8557
rect 22005 8517 22017 8551
rect 22051 8548 22063 8551
rect 22462 8548 22468 8560
rect 22051 8520 22468 8548
rect 22051 8517 22063 8520
rect 22005 8511 22063 8517
rect 22462 8508 22468 8520
rect 22520 8548 22526 8560
rect 22830 8548 22836 8560
rect 22520 8520 22836 8548
rect 22520 8508 22526 8520
rect 22830 8508 22836 8520
rect 22888 8508 22894 8560
rect 23658 8548 23664 8560
rect 23492 8520 23664 8548
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20438 8480 20444 8492
rect 20036 8452 20444 8480
rect 20036 8440 20042 8452
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 20640 8452 21097 8480
rect 13596 8384 14771 8412
rect 15381 8415 15439 8421
rect 13596 8372 13602 8384
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 16666 8412 16672 8424
rect 15427 8384 16672 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 13814 8344 13820 8356
rect 11440 8316 12664 8344
rect 9769 8307 9827 8313
rect 12636 8288 12664 8316
rect 13004 8316 13820 8344
rect 13004 8288 13032 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14826 8344 14832 8356
rect 14787 8316 14832 8344
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 15749 8347 15807 8353
rect 15749 8344 15761 8347
rect 15068 8316 15761 8344
rect 15068 8304 15074 8316
rect 15749 8313 15761 8316
rect 15795 8313 15807 8347
rect 15749 8307 15807 8313
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 17236 8344 17264 8375
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 19245 8415 19303 8421
rect 19245 8412 19257 8415
rect 17920 8384 19257 8412
rect 17920 8372 17926 8384
rect 19245 8381 19257 8384
rect 19291 8381 19303 8415
rect 19245 8375 19303 8381
rect 18046 8344 18052 8356
rect 16356 8316 17172 8344
rect 17236 8316 18052 8344
rect 16356 8304 16362 8316
rect 7340 8248 8524 8276
rect 7340 8236 7346 8248
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 9916 8248 10517 8276
rect 9916 8236 9922 8248
rect 10505 8245 10517 8248
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 12618 8236 12624 8288
rect 12676 8236 12682 8288
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12986 8276 12992 8288
rect 12759 8248 12992 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13449 8279 13507 8285
rect 13449 8276 13461 8279
rect 13320 8248 13461 8276
rect 13320 8236 13326 8248
rect 13449 8245 13461 8248
rect 13495 8245 13507 8279
rect 15562 8276 15568 8288
rect 15523 8248 15568 8276
rect 13449 8239 13507 8245
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16758 8276 16764 8288
rect 16719 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 17144 8276 17172 8316
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 18690 8344 18696 8356
rect 18196 8316 18696 8344
rect 18196 8304 18202 8316
rect 18690 8304 18696 8316
rect 18748 8304 18754 8356
rect 20640 8353 20668 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21416 8452 21833 8480
rect 21416 8440 21422 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22089 8483 22147 8489
rect 22089 8480 22101 8483
rect 21968 8452 22101 8480
rect 21968 8440 21974 8452
rect 22089 8449 22101 8452
rect 22135 8449 22147 8483
rect 22089 8443 22147 8449
rect 22189 8484 22247 8489
rect 22189 8483 22324 8484
rect 22189 8449 22201 8483
rect 22235 8456 22324 8483
rect 22235 8449 22247 8456
rect 22189 8443 22247 8449
rect 22296 8412 22324 8456
rect 22370 8440 22376 8492
rect 22428 8480 22434 8492
rect 23492 8489 23520 8520
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 24762 8548 24768 8560
rect 24596 8520 24768 8548
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22428 8452 23029 8480
rect 22428 8440 22434 8452
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23750 8480 23756 8492
rect 23624 8452 23669 8480
rect 23711 8452 23756 8480
rect 23624 8440 23630 8452
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 23983 8483 24041 8489
rect 23900 8452 23945 8480
rect 23900 8440 23906 8452
rect 23983 8449 23995 8483
rect 24029 8480 24041 8483
rect 24596 8480 24624 8520
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 25884 8548 25912 8588
rect 27246 8576 27252 8588
rect 27304 8576 27310 8628
rect 28166 8576 28172 8628
rect 28224 8616 28230 8628
rect 28224 8588 29316 8616
rect 28224 8576 28230 8588
rect 25756 8520 25912 8548
rect 24029 8452 24624 8480
rect 24029 8449 24041 8452
rect 23983 8443 24041 8449
rect 24670 8440 24676 8492
rect 24728 8480 24734 8492
rect 24728 8452 24773 8480
rect 24728 8440 24734 8452
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25590 8480 25596 8492
rect 25004 8452 25596 8480
rect 25004 8440 25010 8452
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 25756 8489 25784 8520
rect 25958 8508 25964 8560
rect 26016 8548 26022 8560
rect 29017 8551 29075 8557
rect 26016 8520 26061 8548
rect 27540 8520 28304 8548
rect 26016 8508 26022 8520
rect 27540 8492 27568 8520
rect 25741 8483 25799 8489
rect 25741 8449 25753 8483
rect 25787 8449 25799 8483
rect 25741 8443 25799 8449
rect 25869 8483 25927 8489
rect 25869 8449 25881 8483
rect 25915 8449 25927 8483
rect 25869 8443 25927 8449
rect 26099 8483 26157 8489
rect 26099 8449 26111 8483
rect 26145 8480 26157 8483
rect 26602 8480 26608 8492
rect 26145 8452 26608 8480
rect 26145 8449 26157 8452
rect 26099 8443 26157 8449
rect 23106 8412 23112 8424
rect 22296 8384 23112 8412
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 23768 8412 23796 8440
rect 25884 8412 25912 8443
rect 26602 8440 26608 8452
rect 26660 8440 26666 8492
rect 27522 8480 27528 8492
rect 27483 8452 27528 8480
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 27706 8489 27712 8492
rect 27673 8483 27712 8489
rect 27673 8449 27685 8483
rect 27673 8443 27712 8449
rect 27706 8440 27712 8443
rect 27764 8440 27770 8492
rect 27801 8483 27859 8489
rect 27801 8449 27813 8483
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 26694 8412 26700 8424
rect 23768 8384 26700 8412
rect 26694 8372 26700 8384
rect 26752 8372 26758 8424
rect 26786 8372 26792 8424
rect 26844 8412 26850 8424
rect 27816 8412 27844 8443
rect 27890 8440 27896 8492
rect 27948 8480 27954 8492
rect 28031 8483 28089 8489
rect 27948 8452 27993 8480
rect 27948 8440 27954 8452
rect 28031 8449 28043 8483
rect 28077 8480 28089 8483
rect 28166 8480 28172 8492
rect 28077 8452 28172 8480
rect 28077 8449 28089 8452
rect 28031 8443 28089 8449
rect 28166 8440 28172 8452
rect 28224 8440 28230 8492
rect 28276 8480 28304 8520
rect 29017 8517 29029 8551
rect 29063 8548 29075 8551
rect 29178 8548 29184 8560
rect 29063 8520 29184 8548
rect 29063 8517 29075 8520
rect 29017 8511 29075 8517
rect 29178 8508 29184 8520
rect 29236 8508 29242 8560
rect 28810 8489 28816 8492
rect 28618 8483 28676 8489
rect 28276 8478 28488 8480
rect 28618 8478 28630 8483
rect 28276 8452 28630 8478
rect 28460 8450 28630 8452
rect 28618 8449 28630 8450
rect 28664 8449 28676 8483
rect 28618 8443 28676 8449
rect 28777 8483 28816 8489
rect 28777 8449 28789 8483
rect 28777 8443 28816 8449
rect 28810 8440 28816 8443
rect 28868 8440 28874 8492
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29094 8483 29152 8489
rect 28960 8452 29005 8480
rect 28960 8440 28966 8452
rect 29094 8449 29106 8483
rect 29140 8480 29152 8483
rect 29288 8480 29316 8588
rect 30006 8576 30012 8628
rect 30064 8616 30070 8628
rect 30469 8619 30527 8625
rect 30469 8616 30481 8619
rect 30064 8588 30481 8616
rect 30064 8576 30070 8588
rect 30469 8585 30481 8588
rect 30515 8585 30527 8619
rect 30469 8579 30527 8585
rect 30834 8576 30840 8628
rect 30892 8616 30898 8628
rect 34247 8619 34305 8625
rect 30892 8588 33916 8616
rect 30892 8576 30898 8588
rect 32217 8551 32275 8557
rect 32217 8517 32229 8551
rect 32263 8548 32275 8551
rect 32674 8548 32680 8560
rect 32263 8520 32680 8548
rect 32263 8517 32275 8520
rect 32217 8511 32275 8517
rect 32674 8508 32680 8520
rect 32732 8508 32738 8560
rect 33226 8548 33232 8560
rect 33060 8520 33232 8548
rect 30466 8480 30472 8492
rect 29140 8452 29316 8480
rect 30427 8452 30472 8480
rect 29140 8449 29152 8452
rect 29094 8443 29152 8449
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 30837 8483 30895 8489
rect 30837 8449 30849 8483
rect 30883 8480 30895 8483
rect 31110 8480 31116 8492
rect 30883 8452 31116 8480
rect 30883 8449 30895 8452
rect 30837 8443 30895 8449
rect 31110 8440 31116 8452
rect 31168 8440 31174 8492
rect 31386 8480 31392 8492
rect 31347 8452 31392 8480
rect 31386 8440 31392 8452
rect 31444 8440 31450 8492
rect 31478 8440 31484 8492
rect 31536 8480 31542 8492
rect 31573 8483 31631 8489
rect 31573 8480 31585 8483
rect 31536 8452 31585 8480
rect 31536 8440 31542 8452
rect 31573 8449 31585 8452
rect 31619 8449 31631 8483
rect 31573 8443 31631 8449
rect 30558 8412 30564 8424
rect 26844 8384 27844 8412
rect 28966 8384 30564 8412
rect 26844 8372 26850 8384
rect 20625 8347 20683 8353
rect 20625 8313 20637 8347
rect 20671 8313 20683 8347
rect 22370 8344 22376 8356
rect 22331 8316 22376 8344
rect 20625 8307 20683 8313
rect 22370 8304 22376 8316
rect 22428 8344 22434 8356
rect 22646 8344 22652 8356
rect 22428 8316 22652 8344
rect 22428 8304 22434 8316
rect 22646 8304 22652 8316
rect 22704 8304 22710 8356
rect 22830 8344 22836 8356
rect 22791 8316 22836 8344
rect 22830 8304 22836 8316
rect 22888 8304 22894 8356
rect 23124 8344 23152 8372
rect 28966 8356 28994 8384
rect 30558 8372 30564 8384
rect 30616 8372 30622 8424
rect 30742 8372 30748 8424
rect 30800 8412 30806 8424
rect 30929 8415 30987 8421
rect 30929 8412 30941 8415
rect 30800 8384 30941 8412
rect 30800 8372 30806 8384
rect 30929 8381 30941 8384
rect 30975 8381 30987 8415
rect 30929 8375 30987 8381
rect 32677 8415 32735 8421
rect 32677 8381 32689 8415
rect 32723 8412 32735 8415
rect 33060 8412 33088 8520
rect 33226 8508 33232 8520
rect 33284 8508 33290 8560
rect 33502 8508 33508 8560
rect 33560 8508 33566 8560
rect 33134 8440 33140 8492
rect 33192 8480 33198 8492
rect 33321 8483 33379 8489
rect 33192 8452 33272 8480
rect 33192 8440 33198 8452
rect 32723 8384 33088 8412
rect 33244 8412 33272 8452
rect 33321 8449 33333 8483
rect 33367 8480 33379 8483
rect 33520 8480 33548 8508
rect 33367 8452 33548 8480
rect 33367 8449 33379 8452
rect 33321 8443 33379 8449
rect 33413 8415 33471 8421
rect 33413 8412 33425 8415
rect 33244 8384 33425 8412
rect 32723 8381 32735 8384
rect 32677 8375 32735 8381
rect 33413 8381 33425 8384
rect 33459 8381 33471 8415
rect 33413 8375 33471 8381
rect 33505 8415 33563 8421
rect 33505 8381 33517 8415
rect 33551 8381 33563 8415
rect 33505 8375 33563 8381
rect 24854 8344 24860 8356
rect 23124 8316 24860 8344
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 25498 8304 25504 8356
rect 25556 8344 25562 8356
rect 26237 8347 26295 8353
rect 26237 8344 26249 8347
rect 25556 8316 26249 8344
rect 25556 8304 25562 8316
rect 26237 8313 26249 8316
rect 26283 8313 26295 8347
rect 26237 8307 26295 8313
rect 27982 8304 27988 8356
rect 28040 8344 28046 8356
rect 28169 8347 28227 8353
rect 28169 8344 28181 8347
rect 28040 8316 28181 8344
rect 28040 8304 28046 8316
rect 28169 8313 28181 8316
rect 28215 8313 28227 8347
rect 28169 8307 28227 8313
rect 28948 8304 28954 8356
rect 29006 8304 29012 8356
rect 29270 8344 29276 8356
rect 29231 8316 29276 8344
rect 29270 8304 29276 8316
rect 29328 8304 29334 8356
rect 29362 8304 29368 8356
rect 29420 8344 29426 8356
rect 31389 8347 31447 8353
rect 31389 8344 31401 8347
rect 29420 8316 31401 8344
rect 29420 8304 29426 8316
rect 31389 8313 31401 8316
rect 31435 8313 31447 8347
rect 31389 8307 31447 8313
rect 32585 8347 32643 8353
rect 32585 8313 32597 8347
rect 32631 8344 32643 8347
rect 33137 8347 33195 8353
rect 33137 8344 33149 8347
rect 32631 8316 33149 8344
rect 32631 8313 32643 8316
rect 32585 8307 32643 8313
rect 33137 8313 33149 8316
rect 33183 8313 33195 8347
rect 33137 8307 33195 8313
rect 33318 8304 33324 8356
rect 33376 8344 33382 8356
rect 33520 8344 33548 8375
rect 33594 8372 33600 8424
rect 33652 8412 33658 8424
rect 33888 8412 33916 8588
rect 34247 8585 34259 8619
rect 34293 8616 34305 8619
rect 34422 8616 34428 8628
rect 34293 8588 34428 8616
rect 34293 8585 34305 8588
rect 34247 8579 34305 8585
rect 34422 8576 34428 8588
rect 34480 8576 34486 8628
rect 34146 8548 34152 8560
rect 34107 8520 34152 8548
rect 34146 8508 34152 8520
rect 34204 8508 34210 8560
rect 34333 8551 34391 8557
rect 34333 8517 34345 8551
rect 34379 8548 34391 8551
rect 34977 8551 35035 8557
rect 34977 8548 34989 8551
rect 34379 8520 34989 8548
rect 34379 8517 34391 8520
rect 34333 8511 34391 8517
rect 34977 8517 34989 8520
rect 35023 8517 35035 8551
rect 34977 8511 35035 8517
rect 34425 8483 34483 8489
rect 34425 8449 34437 8483
rect 34471 8480 34483 8483
rect 34514 8480 34520 8492
rect 34471 8452 34520 8480
rect 34471 8449 34483 8452
rect 34425 8443 34483 8449
rect 34514 8440 34520 8452
rect 34572 8440 34578 8492
rect 34790 8440 34796 8492
rect 34848 8480 34854 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34848 8452 34897 8480
rect 34848 8440 34854 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 35713 8483 35771 8489
rect 35713 8449 35725 8483
rect 35759 8480 35771 8483
rect 35802 8480 35808 8492
rect 35759 8452 35808 8480
rect 35759 8449 35771 8452
rect 35713 8443 35771 8449
rect 35802 8440 35808 8452
rect 35860 8440 35866 8492
rect 35986 8412 35992 8424
rect 33652 8384 33745 8412
rect 33888 8384 35992 8412
rect 33652 8372 33658 8384
rect 35986 8372 35992 8384
rect 36044 8372 36050 8424
rect 33376 8316 33548 8344
rect 33612 8344 33640 8372
rect 33962 8344 33968 8356
rect 33612 8316 33968 8344
rect 33376 8304 33382 8316
rect 17218 8276 17224 8288
rect 17144 8248 17224 8276
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 18598 8276 18604 8288
rect 18559 8248 18604 8276
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 25590 8236 25596 8288
rect 25648 8276 25654 8288
rect 30006 8276 30012 8288
rect 25648 8248 30012 8276
rect 25648 8236 25654 8248
rect 30006 8236 30012 8248
rect 30064 8236 30070 8288
rect 30285 8279 30343 8285
rect 30285 8245 30297 8279
rect 30331 8276 30343 8279
rect 30374 8276 30380 8288
rect 30331 8248 30380 8276
rect 30331 8245 30343 8248
rect 30285 8239 30343 8245
rect 30374 8236 30380 8248
rect 30432 8236 30438 8288
rect 32306 8236 32312 8288
rect 32364 8276 32370 8288
rect 33410 8276 33416 8288
rect 32364 8248 33416 8276
rect 32364 8236 32370 8248
rect 33410 8236 33416 8248
rect 33468 8236 33474 8288
rect 33520 8276 33548 8316
rect 33962 8304 33968 8316
rect 34020 8304 34026 8356
rect 35618 8344 35624 8356
rect 34072 8316 35624 8344
rect 34072 8276 34100 8316
rect 35618 8304 35624 8316
rect 35676 8304 35682 8356
rect 35526 8276 35532 8288
rect 33520 8248 34100 8276
rect 35487 8248 35532 8276
rect 35526 8236 35532 8248
rect 35584 8236 35590 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 7006 8072 7012 8084
rect 6656 8044 7012 8072
rect 6656 7945 6684 8044
rect 7006 8032 7012 8044
rect 7064 8072 7070 8084
rect 8018 8072 8024 8084
rect 7064 8044 7696 8072
rect 7979 8044 8024 8072
rect 7064 8032 7070 8044
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 7668 7936 7696 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8846 8072 8852 8084
rect 8128 8044 8852 8072
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 8128 8004 8156 8044
rect 8846 8032 8852 8044
rect 8904 8072 8910 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 8904 8044 13369 8072
rect 8904 8032 8910 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 15102 8072 15108 8084
rect 13357 8035 13415 8041
rect 14016 8044 15108 8072
rect 7800 7976 8156 8004
rect 7800 7964 7806 7976
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 7668 7908 9229 7936
rect 6641 7899 6699 7905
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5258 7868 5264 7880
rect 5215 7840 5264 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 6178 7868 6184 7880
rect 5408 7840 5453 7868
rect 6139 7840 6184 7868
rect 5408 7828 5414 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 9232 7868 9260 7899
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 9232 7840 11345 7868
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 14016 7868 14044 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15562 8072 15568 8084
rect 15436 8044 15568 8072
rect 15436 8032 15442 8044
rect 15562 8032 15568 8044
rect 15620 8072 15626 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 15620 8044 17325 8072
rect 15620 8032 15626 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17954 8072 17960 8084
rect 17915 8044 17960 8072
rect 17313 8035 17371 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18414 8072 18420 8084
rect 18279 8044 18420 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 18932 8044 19349 8072
rect 18932 8032 18938 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 23842 8072 23848 8084
rect 23803 8044 23848 8072
rect 19337 8035 19395 8041
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 24762 8072 24768 8084
rect 24627 8044 24768 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 25774 8032 25780 8084
rect 25832 8072 25838 8084
rect 25869 8075 25927 8081
rect 25869 8072 25881 8075
rect 25832 8044 25881 8072
rect 25832 8032 25838 8044
rect 25869 8041 25881 8044
rect 25915 8041 25927 8075
rect 25869 8035 25927 8041
rect 26326 8032 26332 8084
rect 26384 8072 26390 8084
rect 26513 8075 26571 8081
rect 26513 8072 26525 8075
rect 26384 8044 26525 8072
rect 26384 8032 26390 8044
rect 26513 8041 26525 8044
rect 26559 8041 26571 8075
rect 26513 8035 26571 8041
rect 26602 8032 26608 8084
rect 26660 8072 26666 8084
rect 28258 8072 28264 8084
rect 26660 8044 28264 8072
rect 26660 8032 26666 8044
rect 28258 8032 28264 8044
rect 28316 8032 28322 8084
rect 28442 8072 28448 8084
rect 28403 8044 28448 8072
rect 28442 8032 28448 8044
rect 28500 8032 28506 8084
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 30926 8072 30932 8084
rect 28592 8044 30932 8072
rect 28592 8032 28598 8044
rect 30926 8032 30932 8044
rect 30984 8032 30990 8084
rect 31202 8032 31208 8084
rect 31260 8072 31266 8084
rect 31386 8072 31392 8084
rect 31260 8044 31392 8072
rect 31260 8032 31266 8044
rect 31386 8032 31392 8044
rect 31444 8072 31450 8084
rect 35342 8072 35348 8084
rect 31444 8044 35348 8072
rect 31444 8032 31450 8044
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 28166 8004 28172 8016
rect 27264 7976 28172 8004
rect 18598 7936 18604 7948
rect 16960 7908 18604 7936
rect 11333 7831 11391 7837
rect 11440 7840 14044 7868
rect 14093 7871 14151 7877
rect 6908 7803 6966 7809
rect 6908 7769 6920 7803
rect 6954 7800 6966 7803
rect 7190 7800 7196 7812
rect 6954 7772 7196 7800
rect 6954 7769 6966 7772
rect 6908 7763 6966 7769
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 9462 7803 9520 7809
rect 9462 7800 9474 7803
rect 7760 7772 9474 7800
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 7760 7732 7788 7772
rect 9462 7769 9474 7772
rect 9508 7769 9520 7803
rect 11440 7800 11468 7840
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 15930 7868 15936 7880
rect 14139 7840 15936 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16960 7868 16988 7908
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 21818 7936 21824 7948
rect 18748 7908 20116 7936
rect 18748 7896 18754 7908
rect 16132 7840 16988 7868
rect 17773 7871 17831 7877
rect 9462 7763 9520 7769
rect 9646 7772 11468 7800
rect 11600 7803 11658 7809
rect 6043 7704 7788 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 9646 7732 9674 7772
rect 11600 7769 11612 7803
rect 11646 7800 11658 7803
rect 13170 7800 13176 7812
rect 11646 7772 13176 7800
rect 11646 7769 11658 7772
rect 11600 7763 11658 7769
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7769 13323 7803
rect 13265 7763 13323 7769
rect 14360 7803 14418 7809
rect 14360 7769 14372 7803
rect 14406 7800 14418 7803
rect 16132 7800 16160 7840
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 17819 7840 18000 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 14406 7772 16160 7800
rect 16200 7803 16258 7809
rect 14406 7769 14418 7772
rect 14360 7763 14418 7769
rect 16200 7769 16212 7803
rect 16246 7800 16258 7803
rect 17862 7800 17868 7812
rect 16246 7772 17868 7800
rect 16246 7769 16258 7772
rect 16200 7763 16258 7769
rect 8536 7704 9674 7732
rect 8536 7692 8542 7704
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10502 7732 10508 7744
rect 10100 7704 10508 7732
rect 10100 7692 10106 7704
rect 10502 7692 10508 7704
rect 10560 7732 10566 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10560 7704 10609 7732
rect 10560 7692 10566 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12492 7704 12725 7732
rect 12492 7692 12498 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 13280 7732 13308 7763
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 17972 7800 18000 7840
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 20088 7877 20116 7908
rect 21192 7908 21824 7936
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19116 7840 19257 7868
rect 19116 7828 19122 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20990 7868 20996 7880
rect 20073 7831 20131 7837
rect 20180 7840 20996 7868
rect 18046 7800 18052 7812
rect 17972 7772 18052 7800
rect 18046 7760 18052 7772
rect 18104 7800 18110 7812
rect 19444 7800 19472 7831
rect 18104 7772 19472 7800
rect 18104 7760 18110 7772
rect 13354 7732 13360 7744
rect 13267 7704 13360 7732
rect 12713 7695 12771 7701
rect 13354 7692 13360 7704
rect 13412 7732 13418 7744
rect 15102 7732 15108 7744
rect 13412 7704 15108 7732
rect 13412 7692 13418 7704
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 15470 7732 15476 7744
rect 15431 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 20180 7732 20208 7840
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 21192 7877 21220 7908
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 25314 7896 25320 7948
rect 25372 7936 25378 7948
rect 27264 7945 27292 7976
rect 28166 7964 28172 7976
rect 28224 8004 28230 8016
rect 28718 8004 28724 8016
rect 28224 7976 28724 8004
rect 28224 7964 28230 7976
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 30006 8004 30012 8016
rect 29967 7976 30012 8004
rect 30006 7964 30012 7976
rect 30064 7964 30070 8016
rect 32582 8004 32588 8016
rect 30576 7976 32588 8004
rect 27249 7939 27307 7945
rect 25372 7908 25728 7936
rect 25372 7896 25378 7908
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22465 7871 22523 7877
rect 21324 7840 21588 7868
rect 21324 7828 21330 7840
rect 21560 7812 21588 7840
rect 22465 7837 22477 7871
rect 22511 7868 22523 7871
rect 23658 7868 23664 7880
rect 22511 7840 23664 7868
rect 22511 7837 22523 7840
rect 22465 7831 22523 7837
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23808 7840 24409 7868
rect 23808 7828 23814 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 25498 7868 25504 7880
rect 25459 7840 25504 7868
rect 24397 7831 24455 7837
rect 25498 7828 25504 7840
rect 25556 7828 25562 7880
rect 25700 7877 25728 7908
rect 27249 7905 27261 7939
rect 27295 7905 27307 7939
rect 27249 7899 27307 7905
rect 28077 7939 28135 7945
rect 28077 7905 28089 7939
rect 28123 7936 28135 7939
rect 28442 7936 28448 7948
rect 28123 7908 28448 7936
rect 28123 7905 28135 7908
rect 28077 7899 28135 7905
rect 28442 7896 28448 7908
rect 28500 7896 28506 7948
rect 28810 7896 28816 7948
rect 28868 7936 28874 7948
rect 28868 7908 30052 7936
rect 28868 7896 28874 7908
rect 25685 7871 25743 7877
rect 25685 7837 25697 7871
rect 25731 7837 25743 7871
rect 27430 7868 27436 7880
rect 27391 7840 27436 7868
rect 25685 7831 25743 7837
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7837 28319 7871
rect 28261 7831 28319 7837
rect 21542 7760 21548 7812
rect 21600 7800 21606 7812
rect 21637 7803 21695 7809
rect 21637 7800 21649 7803
rect 21600 7772 21649 7800
rect 21600 7760 21606 7772
rect 21637 7769 21649 7772
rect 21683 7769 21695 7803
rect 21637 7763 21695 7769
rect 21726 7760 21732 7812
rect 21784 7800 21790 7812
rect 21821 7803 21879 7809
rect 21821 7800 21833 7803
rect 21784 7772 21833 7800
rect 21784 7760 21790 7772
rect 21821 7769 21833 7772
rect 21867 7769 21879 7803
rect 21821 7763 21879 7769
rect 21910 7760 21916 7812
rect 21968 7800 21974 7812
rect 22710 7803 22768 7809
rect 22710 7800 22722 7803
rect 21968 7772 22722 7800
rect 21968 7760 21974 7772
rect 22710 7769 22722 7772
rect 22756 7769 22768 7803
rect 22710 7763 22768 7769
rect 24670 7760 24676 7812
rect 24728 7800 24734 7812
rect 26421 7803 26479 7809
rect 26421 7800 26433 7803
rect 24728 7772 26433 7800
rect 24728 7760 24734 7772
rect 26421 7769 26433 7772
rect 26467 7769 26479 7803
rect 27448 7800 27476 7828
rect 28276 7800 28304 7831
rect 28350 7828 28356 7880
rect 28408 7868 28414 7880
rect 29825 7871 29883 7877
rect 29825 7868 29837 7871
rect 28408 7840 29837 7868
rect 28408 7828 28414 7840
rect 29825 7837 29837 7840
rect 29871 7837 29883 7871
rect 29825 7831 29883 7837
rect 27448 7772 28304 7800
rect 26421 7763 26479 7769
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 29270 7800 29276 7812
rect 28500 7772 29276 7800
rect 28500 7760 28506 7772
rect 29270 7760 29276 7772
rect 29328 7760 29334 7812
rect 18288 7704 20208 7732
rect 20257 7735 20315 7741
rect 18288 7692 18294 7704
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 20530 7732 20536 7744
rect 20303 7704 20536 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 21174 7732 21180 7744
rect 21135 7704 21180 7732
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 22005 7735 22063 7741
rect 22005 7732 22017 7735
rect 21324 7704 22017 7732
rect 21324 7692 21330 7704
rect 22005 7701 22017 7704
rect 22051 7701 22063 7735
rect 22005 7695 22063 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 24118 7732 24124 7744
rect 23440 7704 24124 7732
rect 23440 7692 23446 7704
rect 24118 7692 24124 7704
rect 24176 7732 24182 7744
rect 27522 7732 27528 7744
rect 24176 7704 27528 7732
rect 24176 7692 24182 7704
rect 27522 7692 27528 7704
rect 27580 7692 27586 7744
rect 27617 7735 27675 7741
rect 27617 7701 27629 7735
rect 27663 7732 27675 7735
rect 28534 7732 28540 7744
rect 27663 7704 28540 7732
rect 27663 7701 27675 7704
rect 27617 7695 27675 7701
rect 28534 7692 28540 7704
rect 28592 7692 28598 7744
rect 29840 7732 29868 7831
rect 30024 7800 30052 7908
rect 30576 7877 30604 7976
rect 32582 7964 32588 7976
rect 32640 7964 32646 8016
rect 30742 7896 30748 7948
rect 30800 7936 30806 7948
rect 30800 7908 31248 7936
rect 30800 7896 30806 7908
rect 30561 7871 30619 7877
rect 30561 7837 30573 7871
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 30650 7828 30656 7880
rect 30708 7868 30714 7880
rect 30926 7868 30932 7880
rect 30708 7840 30753 7868
rect 30887 7840 30932 7868
rect 30708 7828 30714 7840
rect 30926 7828 30932 7840
rect 30984 7828 30990 7880
rect 31110 7868 31116 7880
rect 31071 7840 31116 7868
rect 31110 7828 31116 7840
rect 31168 7828 31174 7880
rect 31220 7868 31248 7908
rect 31570 7896 31576 7948
rect 31628 7936 31634 7948
rect 32309 7939 32367 7945
rect 32309 7936 32321 7939
rect 31628 7908 32321 7936
rect 31628 7896 31634 7908
rect 32309 7905 32321 7908
rect 32355 7936 32367 7939
rect 32490 7936 32496 7948
rect 32355 7908 32496 7936
rect 32355 7905 32367 7908
rect 32309 7899 32367 7905
rect 32490 7896 32496 7908
rect 32548 7896 32554 7948
rect 34054 7896 34060 7948
rect 34112 7936 34118 7948
rect 34112 7908 35572 7936
rect 34112 7896 34118 7908
rect 32033 7871 32091 7877
rect 32033 7868 32045 7871
rect 31220 7840 32045 7868
rect 32033 7837 32045 7840
rect 32079 7837 32091 7871
rect 32033 7831 32091 7837
rect 32122 7828 32128 7880
rect 32180 7868 32186 7880
rect 32398 7868 32404 7880
rect 32180 7840 32225 7868
rect 32359 7840 32404 7868
rect 32180 7828 32186 7840
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 33226 7828 33232 7880
rect 33284 7868 33290 7880
rect 33781 7871 33839 7877
rect 33781 7868 33793 7871
rect 33284 7840 33793 7868
rect 33284 7828 33290 7840
rect 33781 7837 33793 7840
rect 33827 7837 33839 7871
rect 33781 7831 33839 7837
rect 34606 7828 34612 7880
rect 34664 7868 34670 7880
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 34664 7840 34897 7868
rect 34664 7828 34670 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 35342 7868 35348 7880
rect 35303 7840 35348 7868
rect 34885 7831 34943 7837
rect 35342 7828 35348 7840
rect 35400 7828 35406 7880
rect 35544 7877 35572 7908
rect 35529 7871 35587 7877
rect 35529 7837 35541 7871
rect 35575 7837 35587 7871
rect 36170 7868 36176 7880
rect 36131 7840 36176 7868
rect 35529 7831 35587 7837
rect 36170 7828 36176 7840
rect 36228 7828 36234 7880
rect 30668 7800 30696 7828
rect 30834 7800 30840 7812
rect 30024 7772 30696 7800
rect 30795 7772 30840 7800
rect 30834 7760 30840 7772
rect 30892 7760 30898 7812
rect 31018 7760 31024 7812
rect 31076 7800 31082 7812
rect 32953 7803 33011 7809
rect 32953 7800 32965 7803
rect 31076 7772 32965 7800
rect 31076 7760 31082 7772
rect 32953 7769 32965 7772
rect 32999 7769 33011 7803
rect 32953 7763 33011 7769
rect 33410 7760 33416 7812
rect 33468 7800 33474 7812
rect 35437 7803 35495 7809
rect 35437 7800 35449 7803
rect 33468 7772 35449 7800
rect 33468 7760 33474 7772
rect 35437 7769 35449 7772
rect 35483 7769 35495 7803
rect 35437 7763 35495 7769
rect 31386 7732 31392 7744
rect 29840 7704 31392 7732
rect 31386 7692 31392 7704
rect 31444 7692 31450 7744
rect 31849 7735 31907 7741
rect 31849 7701 31861 7735
rect 31895 7732 31907 7735
rect 32030 7732 32036 7744
rect 31895 7704 32036 7732
rect 31895 7701 31907 7704
rect 31849 7695 31907 7701
rect 32030 7692 32036 7704
rect 32088 7692 32094 7744
rect 33042 7732 33048 7744
rect 33003 7704 33048 7732
rect 33042 7692 33048 7704
rect 33100 7692 33106 7744
rect 33594 7732 33600 7744
rect 33555 7704 33600 7732
rect 33594 7692 33600 7704
rect 33652 7692 33658 7744
rect 34514 7692 34520 7744
rect 34572 7732 34578 7744
rect 34701 7735 34759 7741
rect 34701 7732 34713 7735
rect 34572 7704 34713 7732
rect 34572 7692 34578 7704
rect 34701 7701 34713 7704
rect 34747 7701 34759 7735
rect 34701 7695 34759 7701
rect 35710 7692 35716 7744
rect 35768 7732 35774 7744
rect 35989 7735 36047 7741
rect 35989 7732 36001 7735
rect 35768 7704 36001 7732
rect 35768 7692 35774 7704
rect 35989 7701 36001 7704
rect 36035 7701 36047 7735
rect 35989 7695 36047 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 8202 7528 8208 7540
rect 6236 7500 8208 7528
rect 6236 7488 6242 7500
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9582 7528 9588 7540
rect 9171 7500 9588 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9950 7528 9956 7540
rect 9784 7500 9956 7528
rect 5445 7463 5503 7469
rect 5445 7429 5457 7463
rect 5491 7460 5503 7463
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 5491 7432 6561 7460
rect 5491 7429 5503 7432
rect 5445 7423 5503 7429
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 8018 7460 8024 7472
rect 6549 7423 6607 7429
rect 7852 7432 8024 7460
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5408 7364 5641 7392
rect 5408 7352 5414 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 5629 7355 5687 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7101 7395 7159 7401
rect 6880 7364 6925 7392
rect 6880 7352 6886 7364
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7742 7392 7748 7404
rect 7703 7364 7748 7392
rect 7101 7355 7159 7361
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 7116 7324 7144 7355
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 7852 7401 7880 7432
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 8757 7463 8815 7469
rect 8757 7429 8769 7463
rect 8803 7460 8815 7463
rect 9784 7460 9812 7500
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10042 7488 10048 7540
rect 10100 7488 10106 7540
rect 10226 7528 10232 7540
rect 10152 7500 10232 7528
rect 10060 7460 10088 7488
rect 8803 7432 9812 7460
rect 9876 7432 10088 7460
rect 8803 7429 8815 7432
rect 8757 7423 8815 7429
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 8110 7392 8116 7404
rect 8071 7364 8116 7392
rect 7837 7355 7895 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8570 7392 8576 7404
rect 8531 7364 8576 7392
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 9876 7401 9904 7432
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 6052 7296 7144 7324
rect 6052 7284 6058 7296
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 8864 7324 8892 7355
rect 7248 7296 8892 7324
rect 8956 7324 8984 7355
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 10152 7401 10180 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 13538 7528 13544 7540
rect 13499 7500 13544 7528
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14516 7500 15025 7528
rect 14516 7488 14522 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 15102 7488 15108 7540
rect 15160 7488 15166 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 18012 7500 18245 7528
rect 18012 7488 18018 7500
rect 18233 7497 18245 7500
rect 18279 7528 18291 7531
rect 19058 7528 19064 7540
rect 18279 7500 19064 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 21085 7531 21143 7537
rect 19168 7500 21036 7528
rect 12069 7463 12127 7469
rect 12069 7429 12081 7463
rect 12115 7460 12127 7463
rect 12618 7460 12624 7472
rect 12115 7432 12624 7460
rect 12115 7429 12127 7432
rect 12069 7423 12127 7429
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 13173 7463 13231 7469
rect 13173 7429 13185 7463
rect 13219 7460 13231 7463
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 13219 7432 14013 7460
rect 13219 7429 13231 7432
rect 13173 7423 13231 7429
rect 14001 7429 14013 7432
rect 14047 7429 14059 7463
rect 15120 7460 15148 7488
rect 16390 7460 16396 7472
rect 15120 7432 16396 7460
rect 14001 7423 14059 7429
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 10008 7364 10057 7392
rect 10008 7352 10014 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12526 7392 12532 7404
rect 12299 7364 12532 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 10244 7324 10272 7355
rect 12526 7352 12532 7364
rect 12584 7392 12590 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12584 7364 13369 7392
rect 12584 7352 12590 7364
rect 13357 7361 13369 7364
rect 13403 7392 13415 7395
rect 13446 7392 13452 7404
rect 13403 7364 13452 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7392 14611 7395
rect 14918 7392 14924 7404
rect 14599 7364 14924 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 8956 7296 10272 7324
rect 7248 7284 7254 7296
rect 10060 7268 10088 7296
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 13262 7324 13268 7336
rect 12768 7296 13268 7324
rect 12768 7284 12774 7296
rect 13262 7284 13268 7296
rect 13320 7324 13326 7336
rect 14200 7324 14228 7355
rect 13320 7296 14228 7324
rect 14292 7324 14320 7355
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15212 7401 15240 7432
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 16758 7420 16764 7472
rect 16816 7460 16822 7472
rect 17098 7463 17156 7469
rect 17098 7460 17110 7463
rect 16816 7432 17110 7460
rect 16816 7420 16822 7432
rect 17098 7429 17110 7432
rect 17144 7429 17156 7463
rect 17098 7423 17156 7429
rect 15198 7395 15256 7401
rect 15198 7361 15210 7395
rect 15244 7361 15256 7395
rect 15198 7355 15256 7361
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15378 7392 15384 7404
rect 15335 7364 15384 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 15988 7364 16865 7392
rect 15988 7352 15994 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17402 7352 17408 7404
rect 17460 7392 17466 7404
rect 17460 7364 18460 7392
rect 17460 7352 17466 7364
rect 15470 7324 15476 7336
rect 14292 7296 15476 7324
rect 13320 7284 13326 7296
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 18432 7324 18460 7364
rect 18506 7352 18512 7404
rect 18564 7392 18570 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18564 7364 19073 7392
rect 18564 7352 18570 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 18785 7327 18843 7333
rect 18785 7324 18797 7327
rect 18432 7296 18797 7324
rect 18785 7293 18797 7296
rect 18831 7324 18843 7327
rect 19168 7324 19196 7500
rect 19518 7460 19524 7472
rect 19260 7432 19524 7460
rect 19260 7401 19288 7432
rect 19518 7420 19524 7432
rect 19576 7460 19582 7472
rect 20162 7460 20168 7472
rect 19576 7432 20168 7460
rect 19576 7420 19582 7432
rect 20162 7420 20168 7432
rect 20220 7420 20226 7472
rect 20622 7460 20628 7472
rect 20272 7432 20628 7460
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19978 7392 19984 7404
rect 19659 7364 19984 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20272 7401 20300 7432
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 21008 7460 21036 7500
rect 21085 7497 21097 7531
rect 21131 7528 21143 7531
rect 21818 7528 21824 7540
rect 21131 7500 21824 7528
rect 21131 7497 21143 7500
rect 21085 7491 21143 7497
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 22520 7500 24532 7528
rect 22520 7488 22526 7500
rect 23293 7463 23351 7469
rect 23293 7460 23305 7463
rect 21008 7432 21864 7460
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 21266 7392 21272 7404
rect 21227 7364 21272 7392
rect 20441 7355 20499 7361
rect 18831 7296 19196 7324
rect 19521 7327 19579 7333
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 19521 7293 19533 7327
rect 19567 7324 19579 7327
rect 20162 7324 20168 7336
rect 19567 7296 20168 7324
rect 19567 7293 19579 7296
rect 19521 7287 19579 7293
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 7055 7228 8033 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 8021 7225 8033 7228
rect 8067 7256 8079 7259
rect 9858 7256 9864 7268
rect 8067 7228 9864 7256
rect 8067 7225 8079 7228
rect 8021 7219 8079 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10042 7216 10048 7268
rect 10100 7216 10106 7268
rect 12437 7259 12495 7265
rect 12437 7225 12449 7259
rect 12483 7256 12495 7259
rect 14918 7256 14924 7268
rect 12483 7228 14924 7256
rect 12483 7225 12495 7228
rect 12437 7219 12495 7225
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 18874 7256 18880 7268
rect 18835 7228 18880 7256
rect 18874 7216 18880 7228
rect 18932 7256 18938 7268
rect 20456 7256 20484 7355
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21836 7401 21864 7432
rect 22066 7432 23305 7460
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22066 7392 22094 7432
rect 23293 7429 23305 7432
rect 23339 7460 23351 7463
rect 24394 7460 24400 7472
rect 23339 7432 24400 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 21867 7364 22094 7392
rect 22281 7395 22339 7401
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22462 7392 22468 7404
rect 22327 7364 22468 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 22060 7296 22109 7324
rect 22060 7284 22066 7296
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 22738 7284 22744 7336
rect 22796 7324 22802 7336
rect 22848 7324 22876 7355
rect 23382 7352 23388 7404
rect 23440 7392 23446 7404
rect 23477 7395 23535 7401
rect 23477 7392 23489 7395
rect 23440 7364 23489 7392
rect 23440 7352 23446 7364
rect 23477 7361 23489 7364
rect 23523 7361 23535 7395
rect 23477 7355 23535 7361
rect 23569 7395 23627 7401
rect 23569 7361 23581 7395
rect 23615 7392 23627 7395
rect 23934 7392 23940 7404
rect 23615 7364 23940 7392
rect 23615 7361 23627 7364
rect 23569 7355 23627 7361
rect 23934 7352 23940 7364
rect 23992 7352 23998 7404
rect 24504 7392 24532 7500
rect 24854 7488 24860 7540
rect 24912 7528 24918 7540
rect 27338 7528 27344 7540
rect 24912 7500 27344 7528
rect 24912 7488 24918 7500
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28445 7531 28503 7537
rect 28445 7528 28457 7531
rect 27948 7500 28457 7528
rect 27948 7488 27954 7500
rect 28445 7497 28457 7500
rect 28491 7497 28503 7531
rect 28445 7491 28503 7497
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 29052 7500 29101 7528
rect 29052 7488 29058 7500
rect 29089 7497 29101 7500
rect 29135 7528 29147 7531
rect 30742 7528 30748 7540
rect 29135 7500 30748 7528
rect 29135 7497 29147 7500
rect 29089 7491 29147 7497
rect 30742 7488 30748 7500
rect 30800 7488 30806 7540
rect 30926 7488 30932 7540
rect 30984 7528 30990 7540
rect 31205 7531 31263 7537
rect 31205 7528 31217 7531
rect 30984 7500 31217 7528
rect 30984 7488 30990 7500
rect 31205 7497 31217 7500
rect 31251 7497 31263 7531
rect 31205 7491 31263 7497
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 35342 7528 35348 7540
rect 31444 7500 35348 7528
rect 31444 7488 31450 7500
rect 35342 7488 35348 7500
rect 35400 7488 35406 7540
rect 26237 7463 26295 7469
rect 26237 7429 26249 7463
rect 26283 7460 26295 7463
rect 26786 7460 26792 7472
rect 26283 7432 26792 7460
rect 26283 7429 26295 7432
rect 26237 7423 26295 7429
rect 26786 7420 26792 7432
rect 26844 7420 26850 7472
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 31846 7460 31852 7472
rect 27488 7432 28948 7460
rect 27488 7420 27494 7432
rect 24854 7392 24860 7404
rect 24504 7364 24860 7392
rect 24854 7352 24860 7364
rect 24912 7392 24918 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24912 7364 25053 7392
rect 24912 7352 24918 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25590 7392 25596 7404
rect 25551 7364 25596 7392
rect 25409 7355 25467 7361
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 22796 7296 23520 7324
rect 22796 7284 22802 7296
rect 18932 7228 20484 7256
rect 18932 7216 18938 7228
rect 21450 7216 21456 7268
rect 21508 7256 21514 7268
rect 21910 7256 21916 7268
rect 21508 7228 21916 7256
rect 21508 7216 21514 7228
rect 21910 7216 21916 7228
rect 21968 7216 21974 7268
rect 23382 7256 23388 7268
rect 22066 7228 23388 7256
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6546 7188 6552 7200
rect 5859 7160 6552 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 7558 7188 7564 7200
rect 7519 7160 7564 7188
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 9732 7160 10425 7188
rect 9732 7148 9738 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 14366 7188 14372 7200
rect 12860 7160 14372 7188
rect 12860 7148 12866 7160
rect 14366 7148 14372 7160
rect 14424 7188 14430 7200
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14424 7160 14473 7188
rect 14424 7148 14430 7160
rect 14461 7157 14473 7160
rect 14507 7188 14519 7191
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 14507 7160 15485 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 15473 7157 15485 7160
rect 15519 7188 15531 7191
rect 15838 7188 15844 7200
rect 15519 7160 15844 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15838 7148 15844 7160
rect 15896 7188 15902 7200
rect 16206 7188 16212 7200
rect 15896 7160 16212 7188
rect 15896 7148 15902 7160
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20530 7148 20536 7200
rect 20588 7188 20594 7200
rect 22066 7188 22094 7228
rect 23382 7216 23388 7228
rect 23440 7216 23446 7268
rect 23290 7188 23296 7200
rect 20588 7160 22094 7188
rect 23251 7160 23296 7188
rect 20588 7148 20594 7160
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 23492 7188 23520 7296
rect 23584 7296 24593 7324
rect 23584 7268 23612 7296
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 25130 7324 25136 7336
rect 25091 7296 25136 7324
rect 24581 7287 24639 7293
rect 25130 7284 25136 7296
rect 25188 7284 25194 7336
rect 25424 7324 25452 7355
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 28920 7401 28948 7432
rect 29840 7432 31852 7460
rect 29840 7404 29868 7432
rect 31846 7420 31852 7432
rect 31904 7460 31910 7472
rect 33042 7460 33048 7472
rect 31904 7432 33048 7460
rect 31904 7420 31910 7432
rect 27332 7395 27390 7401
rect 27332 7361 27344 7395
rect 27378 7392 27390 7395
rect 28905 7395 28963 7401
rect 27378 7364 28856 7392
rect 27378 7361 27390 7364
rect 27332 7355 27390 7361
rect 26050 7324 26056 7336
rect 25424 7296 26056 7324
rect 26050 7284 26056 7296
rect 26108 7284 26114 7336
rect 27062 7324 27068 7336
rect 27023 7296 27068 7324
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 23566 7216 23572 7268
rect 23624 7216 23630 7268
rect 24673 7259 24731 7265
rect 24673 7225 24685 7259
rect 24719 7256 24731 7259
rect 26421 7259 26479 7265
rect 24719 7228 26372 7256
rect 24719 7225 24731 7228
rect 24673 7219 24731 7225
rect 25590 7188 25596 7200
rect 23492 7160 25596 7188
rect 25590 7148 25596 7160
rect 25648 7148 25654 7200
rect 26344 7188 26372 7228
rect 26421 7225 26433 7259
rect 26467 7256 26479 7259
rect 26786 7256 26792 7268
rect 26467 7228 26792 7256
rect 26467 7225 26479 7228
rect 26421 7219 26479 7225
rect 26786 7216 26792 7228
rect 26844 7216 26850 7268
rect 28828 7256 28856 7364
rect 28905 7361 28917 7395
rect 28951 7361 28963 7395
rect 29822 7392 29828 7404
rect 29735 7364 29828 7392
rect 28905 7355 28963 7361
rect 29822 7352 29828 7364
rect 29880 7352 29886 7404
rect 30092 7395 30150 7401
rect 30092 7361 30104 7395
rect 30138 7392 30150 7395
rect 32306 7392 32312 7404
rect 30138 7364 32312 7392
rect 30138 7361 30150 7364
rect 30092 7355 30150 7361
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 32600 7401 32628 7432
rect 33042 7420 33048 7432
rect 33100 7460 33106 7472
rect 34968 7463 35026 7469
rect 33100 7432 34744 7460
rect 33100 7420 33106 7432
rect 34716 7404 34744 7432
rect 34968 7429 34980 7463
rect 35014 7460 35026 7463
rect 35526 7460 35532 7472
rect 35014 7432 35532 7460
rect 35014 7429 35026 7432
rect 34968 7423 35026 7429
rect 35526 7420 35532 7432
rect 35584 7420 35590 7472
rect 32585 7395 32643 7401
rect 32585 7361 32597 7395
rect 32631 7361 32643 7395
rect 32585 7355 32643 7361
rect 32852 7395 32910 7401
rect 32852 7361 32864 7395
rect 32898 7392 32910 7395
rect 33594 7392 33600 7404
rect 32898 7364 33600 7392
rect 32898 7361 32910 7364
rect 32852 7355 32910 7361
rect 33594 7352 33600 7364
rect 33652 7352 33658 7404
rect 34698 7392 34704 7404
rect 34611 7364 34704 7392
rect 34698 7352 34704 7364
rect 34756 7352 34762 7404
rect 28828 7228 29592 7256
rect 28626 7188 28632 7200
rect 26344 7160 28632 7188
rect 28626 7148 28632 7160
rect 28684 7148 28690 7200
rect 29564 7188 29592 7228
rect 33888 7228 34744 7256
rect 33888 7188 33916 7228
rect 29564 7160 33916 7188
rect 33962 7148 33968 7200
rect 34020 7188 34026 7200
rect 34716 7188 34744 7228
rect 35894 7188 35900 7200
rect 34020 7160 34065 7188
rect 34716 7160 35900 7188
rect 34020 7148 34026 7160
rect 35894 7148 35900 7160
rect 35952 7148 35958 7200
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 36081 7191 36139 7197
rect 36081 7188 36093 7191
rect 36044 7160 36093 7188
rect 36044 7148 36050 7160
rect 36081 7157 36093 7160
rect 36127 7157 36139 7191
rect 36081 7151 36139 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 6641 6987 6699 6993
rect 5224 6956 6224 6984
rect 5224 6944 5230 6956
rect 6196 6916 6224 6956
rect 6641 6953 6653 6987
rect 6687 6984 6699 6987
rect 6822 6984 6828 6996
rect 6687 6956 6828 6984
rect 6687 6953 6699 6956
rect 6641 6947 6699 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 17494 6984 17500 6996
rect 13228 6956 17500 6984
rect 13228 6944 13234 6956
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 18414 6984 18420 6996
rect 17972 6956 18420 6984
rect 10226 6916 10232 6928
rect 6196 6888 10232 6916
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 16206 6916 16212 6928
rect 12492 6888 13023 6916
rect 16167 6888 16212 6916
rect 12492 6876 12498 6888
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 4948 6820 5273 6848
rect 4948 6808 4954 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 5261 6811 5319 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 8260 6820 9321 6848
rect 8260 6808 8266 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9766 6848 9772 6860
rect 9727 6820 9772 6848
rect 9309 6811 9367 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 11698 6848 11704 6860
rect 11379 6820 11704 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11698 6808 11704 6820
rect 11756 6848 11762 6860
rect 12342 6848 12348 6860
rect 11756 6820 12348 6848
rect 11756 6808 11762 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12618 6848 12624 6860
rect 12579 6820 12624 6848
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7558 6780 7564 6792
rect 7147 6752 7564 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8662 6780 8668 6792
rect 8343 6752 8668 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9674 6780 9680 6792
rect 9171 6752 9680 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 5528 6715 5586 6721
rect 5528 6681 5540 6715
rect 5574 6712 5586 6715
rect 6362 6712 6368 6724
rect 5574 6684 6368 6712
rect 5574 6681 5586 6684
rect 5528 6675 5586 6681
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 7282 6712 7288 6724
rect 7243 6684 7288 6712
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 9048 6712 9076 6743
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11606 6780 11612 6792
rect 11567 6752 11612 6780
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12995 6789 13023 6888
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 16390 6876 16396 6928
rect 16448 6916 16454 6928
rect 16761 6919 16819 6925
rect 16761 6916 16773 6919
rect 16448 6888 16773 6916
rect 16448 6876 16454 6888
rect 16761 6885 16773 6888
rect 16807 6885 16819 6919
rect 17972 6916 18000 6956
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 21174 6944 21180 6996
rect 21232 6984 21238 6996
rect 21913 6987 21971 6993
rect 21232 6956 21588 6984
rect 21232 6944 21238 6956
rect 19702 6916 19708 6928
rect 16761 6879 16819 6885
rect 17880 6888 18000 6916
rect 18340 6888 19708 6916
rect 13081 6851 13139 6857
rect 13081 6817 13093 6851
rect 13127 6848 13139 6851
rect 13127 6820 13492 6848
rect 13127 6817 13139 6820
rect 13081 6811 13139 6817
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 12768 6752 12817 6780
rect 12768 6740 12774 6752
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12957 6783 13023 6789
rect 12957 6749 12969 6783
rect 13003 6752 13023 6783
rect 13173 6783 13231 6789
rect 13003 6749 13015 6752
rect 12957 6743 13015 6749
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13464 6780 13492 6820
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 14332 6820 15393 6848
rect 14332 6808 14338 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 17880 6848 17908 6888
rect 18046 6848 18052 6860
rect 15381 6811 15439 6817
rect 16868 6820 17908 6848
rect 18007 6820 18052 6848
rect 13814 6780 13820 6792
rect 13464 6752 13820 6780
rect 13173 6743 13231 6749
rect 9398 6712 9404 6724
rect 8076 6684 9404 6712
rect 8076 6672 8082 6684
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 13188 6712 13216 6743
rect 13814 6740 13820 6752
rect 13872 6780 13878 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 13872 6752 14565 6780
rect 13872 6740 13878 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 14553 6743 14611 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6780 16083 6783
rect 16666 6780 16672 6792
rect 16071 6752 16672 6780
rect 16071 6749 16083 6752
rect 16025 6743 16083 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16868 6789 16896 6820
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 17954 6780 17960 6792
rect 17915 6752 17960 6780
rect 16853 6743 16911 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18340 6780 18368 6888
rect 19702 6876 19708 6888
rect 19760 6876 19766 6928
rect 21560 6916 21588 6956
rect 21913 6953 21925 6987
rect 21959 6984 21971 6987
rect 22646 6984 22652 6996
rect 21959 6956 22652 6984
rect 21959 6953 21971 6956
rect 21913 6947 21971 6953
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 22922 6984 22928 6996
rect 22883 6956 22928 6984
rect 22922 6944 22928 6956
rect 22980 6944 22986 6996
rect 23477 6987 23535 6993
rect 23477 6953 23489 6987
rect 23523 6984 23535 6987
rect 23566 6984 23572 6996
rect 23523 6956 23572 6984
rect 23523 6953 23535 6956
rect 23477 6947 23535 6953
rect 23566 6944 23572 6956
rect 23624 6944 23630 6996
rect 26510 6984 26516 6996
rect 24504 6956 26516 6984
rect 21560 6888 22094 6916
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 18472 6820 20545 6848
rect 18472 6808 18478 6820
rect 20533 6817 20545 6820
rect 20579 6817 20591 6851
rect 22066 6848 22094 6888
rect 22554 6876 22560 6928
rect 22612 6916 22618 6928
rect 24504 6925 24532 6956
rect 26510 6944 26516 6956
rect 26568 6944 26574 6996
rect 26789 6987 26847 6993
rect 26789 6953 26801 6987
rect 26835 6984 26847 6987
rect 27430 6984 27436 6996
rect 26835 6956 27436 6984
rect 26835 6953 26847 6956
rect 26789 6947 26847 6953
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 27522 6944 27528 6996
rect 27580 6984 27586 6996
rect 31570 6984 31576 6996
rect 27580 6956 31576 6984
rect 27580 6944 27586 6956
rect 31570 6944 31576 6956
rect 31628 6944 31634 6996
rect 31846 6984 31852 6996
rect 31680 6956 31852 6984
rect 24489 6919 24547 6925
rect 22612 6888 22784 6916
rect 22612 6876 22618 6888
rect 22756 6848 22784 6888
rect 24489 6885 24501 6919
rect 24535 6885 24547 6919
rect 24489 6879 24547 6885
rect 30009 6919 30067 6925
rect 30009 6885 30021 6919
rect 30055 6916 30067 6919
rect 31478 6916 31484 6928
rect 30055 6888 31484 6916
rect 30055 6885 30067 6888
rect 30009 6879 30067 6885
rect 31478 6876 31484 6888
rect 31536 6876 31542 6928
rect 23017 6851 23075 6857
rect 23017 6848 23029 6851
rect 22066 6820 22692 6848
rect 22756 6820 23029 6848
rect 20533 6811 20591 6817
rect 22664 6792 22692 6820
rect 23017 6817 23029 6820
rect 23063 6817 23075 6851
rect 23934 6848 23940 6860
rect 23017 6811 23075 6817
rect 23492 6820 23940 6848
rect 18064 6752 18368 6780
rect 14182 6712 14188 6724
rect 12308 6684 13216 6712
rect 13648 6684 14188 6712
rect 12308 6672 12314 6684
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 7892 6616 8125 6644
rect 7892 6604 7898 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 13648 6644 13676 6684
rect 14182 6672 14188 6684
rect 14240 6672 14246 6724
rect 14366 6712 14372 6724
rect 14327 6684 14372 6712
rect 14366 6672 14372 6684
rect 14424 6672 14430 6724
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15197 6715 15255 6721
rect 15197 6712 15209 6715
rect 15160 6684 15209 6712
rect 15160 6672 15166 6684
rect 15197 6681 15209 6684
rect 15243 6681 15255 6715
rect 18064 6712 18092 6752
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 18748 6752 19441 6780
rect 18748 6740 18754 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 20073 6783 20131 6789
rect 20073 6780 20085 6783
rect 19760 6752 20085 6780
rect 19760 6740 19766 6752
rect 20073 6749 20085 6752
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22498 6783 22556 6789
rect 22498 6780 22510 6783
rect 21968 6752 22510 6780
rect 21968 6740 21974 6752
rect 22498 6749 22510 6752
rect 22544 6749 22556 6783
rect 22498 6743 22556 6749
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 23492 6789 23520 6820
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 24394 6848 24400 6860
rect 24355 6820 24400 6848
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 24578 6808 24584 6860
rect 24636 6848 24642 6860
rect 24765 6851 24823 6857
rect 24765 6848 24777 6851
rect 24636 6820 24777 6848
rect 24636 6808 24642 6820
rect 24765 6817 24777 6820
rect 24811 6817 24823 6851
rect 24765 6811 24823 6817
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 30650 6848 30656 6860
rect 27396 6820 28488 6848
rect 27396 6808 27402 6820
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 24670 6780 24676 6792
rect 23707 6752 24676 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 24854 6780 24860 6792
rect 24815 6752 24860 6780
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 25188 6752 25237 6780
rect 25188 6740 25194 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6780 25467 6783
rect 25590 6780 25596 6792
rect 25455 6752 25596 6780
rect 25455 6749 25467 6752
rect 25409 6743 25467 6749
rect 25590 6740 25596 6752
rect 25648 6740 25654 6792
rect 26326 6780 26332 6792
rect 26287 6752 26332 6780
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 18230 6712 18236 6724
rect 15197 6675 15255 6681
rect 17788 6684 18092 6712
rect 18191 6684 18236 6712
rect 9824 6616 13676 6644
rect 9824 6604 9830 6616
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 14642 6644 14648 6656
rect 13780 6616 14648 6644
rect 13780 6604 13786 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 17788 6644 17816 6684
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 18322 6672 18328 6724
rect 18380 6712 18386 6724
rect 20800 6715 20858 6721
rect 18380 6684 18425 6712
rect 18524 6684 19932 6712
rect 18380 6672 18386 6684
rect 14884 6616 17816 6644
rect 14884 6604 14890 6616
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 18524 6644 18552 6684
rect 19242 6644 19248 6656
rect 17920 6616 18552 6644
rect 19203 6616 19248 6644
rect 17920 6604 17926 6616
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19904 6653 19932 6684
rect 20800 6681 20812 6715
rect 20846 6712 20858 6715
rect 20898 6712 20904 6724
rect 20846 6684 20904 6712
rect 20846 6681 20858 6684
rect 20800 6675 20858 6681
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 23106 6672 23112 6724
rect 23164 6712 23170 6724
rect 26804 6712 26832 6743
rect 26878 6740 26884 6792
rect 26936 6780 26942 6792
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 26936 6752 26985 6780
rect 26936 6740 26942 6752
rect 26973 6749 26985 6752
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 27062 6740 27068 6792
rect 27120 6780 27126 6792
rect 27430 6780 27436 6792
rect 27120 6752 27436 6780
rect 27120 6740 27126 6752
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6780 27859 6783
rect 27890 6780 27896 6792
rect 27847 6752 27896 6780
rect 27847 6749 27859 6752
rect 27801 6743 27859 6749
rect 27890 6740 27896 6752
rect 27948 6740 27954 6792
rect 28460 6789 28488 6820
rect 29932 6820 30656 6848
rect 28445 6783 28503 6789
rect 28445 6749 28457 6783
rect 28491 6780 28503 6783
rect 28534 6780 28540 6792
rect 28491 6752 28540 6780
rect 28491 6749 28503 6752
rect 28445 6743 28503 6749
rect 28534 6740 28540 6752
rect 28592 6740 28598 6792
rect 29730 6780 29736 6792
rect 29691 6752 29736 6780
rect 29730 6740 29736 6752
rect 29788 6740 29794 6792
rect 29932 6789 29960 6820
rect 30650 6808 30656 6820
rect 30708 6808 30714 6860
rect 31202 6848 31208 6860
rect 31163 6820 31208 6848
rect 31202 6808 31208 6820
rect 31260 6808 31266 6860
rect 31680 6857 31708 6956
rect 31846 6944 31852 6956
rect 31904 6984 31910 6996
rect 32306 6984 32312 6996
rect 31904 6956 32312 6984
rect 31904 6944 31910 6956
rect 32306 6944 32312 6956
rect 32364 6944 32370 6996
rect 32398 6944 32404 6996
rect 32456 6984 32462 6996
rect 33045 6987 33103 6993
rect 33045 6984 33057 6987
rect 32456 6956 33057 6984
rect 32456 6944 32462 6956
rect 33045 6953 33057 6956
rect 33091 6953 33103 6987
rect 35710 6984 35716 6996
rect 33045 6947 33103 6953
rect 33152 6956 35716 6984
rect 33152 6916 33180 6956
rect 35710 6944 35716 6956
rect 35768 6944 35774 6996
rect 35894 6984 35900 6996
rect 35855 6956 35900 6984
rect 35894 6944 35900 6956
rect 35952 6944 35958 6996
rect 33060 6888 33180 6916
rect 31665 6851 31723 6857
rect 31665 6817 31677 6851
rect 31711 6817 31723 6851
rect 31665 6811 31723 6817
rect 29917 6783 29975 6789
rect 29917 6749 29929 6783
rect 29963 6749 29975 6783
rect 30190 6780 30196 6792
rect 30151 6752 30196 6780
rect 29917 6743 29975 6749
rect 30190 6740 30196 6752
rect 30248 6740 30254 6792
rect 30466 6780 30472 6792
rect 30427 6752 30472 6780
rect 30466 6740 30472 6752
rect 30524 6740 30530 6792
rect 31932 6783 31990 6789
rect 31932 6749 31944 6783
rect 31978 6780 31990 6783
rect 33060 6780 33088 6888
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 35434 6848 35440 6860
rect 33192 6820 35440 6848
rect 33192 6808 33198 6820
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 31978 6752 33088 6780
rect 33689 6783 33747 6789
rect 31978 6749 31990 6752
rect 31932 6743 31990 6749
rect 33689 6749 33701 6783
rect 33735 6749 33747 6783
rect 33689 6743 33747 6749
rect 27614 6712 27620 6724
rect 23164 6684 26832 6712
rect 27575 6684 27620 6712
rect 23164 6672 23170 6684
rect 27614 6672 27620 6684
rect 27672 6672 27678 6724
rect 27982 6712 27988 6724
rect 27943 6684 27988 6712
rect 27982 6672 27988 6684
rect 28040 6672 28046 6724
rect 28258 6672 28264 6724
rect 28316 6712 28322 6724
rect 31021 6715 31079 6721
rect 31021 6712 31033 6715
rect 28316 6684 31033 6712
rect 28316 6672 28322 6684
rect 31021 6681 31033 6684
rect 31067 6712 31079 6715
rect 33134 6712 33140 6724
rect 31067 6684 33140 6712
rect 31067 6681 31079 6684
rect 31021 6675 31079 6681
rect 33134 6672 33140 6684
rect 33192 6672 33198 6724
rect 33226 6672 33232 6724
rect 33284 6712 33290 6724
rect 33704 6712 33732 6743
rect 34790 6740 34796 6792
rect 34848 6780 34854 6792
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 34848 6752 34897 6780
rect 34848 6740 34854 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 35250 6780 35256 6792
rect 35211 6752 35256 6780
rect 34885 6743 34943 6749
rect 35250 6740 35256 6752
rect 35308 6740 35314 6792
rect 36262 6780 36268 6792
rect 36081 6759 36139 6765
rect 36081 6725 36093 6759
rect 36127 6756 36139 6759
rect 36188 6756 36268 6780
rect 36127 6752 36268 6756
rect 36127 6728 36216 6752
rect 36262 6740 36268 6752
rect 36320 6740 36326 6792
rect 36722 6780 36728 6792
rect 36683 6752 36728 6780
rect 36722 6740 36728 6752
rect 36780 6740 36786 6792
rect 37366 6780 37372 6792
rect 37327 6752 37372 6780
rect 37366 6740 37372 6752
rect 37424 6740 37430 6792
rect 36127 6725 36139 6728
rect 35066 6712 35072 6724
rect 33284 6684 33732 6712
rect 35027 6684 35072 6712
rect 33284 6672 33290 6684
rect 35066 6672 35072 6684
rect 35124 6672 35130 6724
rect 35161 6715 35219 6721
rect 35161 6681 35173 6715
rect 35207 6712 35219 6715
rect 35986 6712 35992 6724
rect 35207 6684 35992 6712
rect 35207 6681 35219 6684
rect 35161 6675 35219 6681
rect 35986 6672 35992 6684
rect 36044 6672 36050 6724
rect 36081 6719 36139 6725
rect 19889 6647 19947 6653
rect 19889 6613 19901 6647
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 22373 6647 22431 6653
rect 22373 6613 22385 6647
rect 22419 6644 22431 6647
rect 22462 6644 22468 6656
rect 22419 6616 22468 6644
rect 22419 6613 22431 6616
rect 22373 6607 22431 6613
rect 22462 6604 22468 6616
rect 22520 6604 22526 6656
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6644 22615 6647
rect 22738 6644 22744 6656
rect 22603 6616 22744 6644
rect 22603 6613 22615 6616
rect 22557 6607 22615 6613
rect 22738 6604 22744 6616
rect 22796 6604 22802 6656
rect 24578 6604 24584 6656
rect 24636 6644 24642 6656
rect 26145 6647 26203 6653
rect 26145 6644 26157 6647
rect 24636 6616 26157 6644
rect 24636 6604 24642 6616
rect 26145 6613 26157 6616
rect 26191 6613 26203 6647
rect 26145 6607 26203 6613
rect 28442 6604 28448 6656
rect 28500 6644 28506 6656
rect 28629 6647 28687 6653
rect 28629 6644 28641 6647
rect 28500 6616 28641 6644
rect 28500 6604 28506 6616
rect 28629 6613 28641 6616
rect 28675 6644 28687 6647
rect 30466 6644 30472 6656
rect 28675 6616 30472 6644
rect 28675 6613 28687 6616
rect 28629 6607 28687 6613
rect 30466 6604 30472 6616
rect 30524 6644 30530 6656
rect 30926 6644 30932 6656
rect 30524 6616 30932 6644
rect 30524 6604 30530 6616
rect 30926 6604 30932 6616
rect 30984 6644 30990 6656
rect 31110 6644 31116 6656
rect 30984 6616 31116 6644
rect 30984 6604 30990 6616
rect 31110 6604 31116 6616
rect 31168 6604 31174 6656
rect 33502 6644 33508 6656
rect 33463 6616 33508 6644
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 35437 6647 35495 6653
rect 35437 6613 35449 6647
rect 35483 6644 35495 6647
rect 35894 6644 35900 6656
rect 35483 6616 35900 6644
rect 35483 6613 35495 6616
rect 35437 6607 35495 6613
rect 35894 6604 35900 6616
rect 35952 6604 35958 6656
rect 36262 6604 36268 6656
rect 36320 6644 36326 6656
rect 36541 6647 36599 6653
rect 36541 6644 36553 6647
rect 36320 6616 36553 6644
rect 36320 6604 36326 6616
rect 36541 6613 36553 6616
rect 36587 6613 36599 6647
rect 37182 6644 37188 6656
rect 37143 6616 37188 6644
rect 36541 6607 36599 6613
rect 37182 6604 37188 6616
rect 37240 6604 37246 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4706 6440 4712 6452
rect 4387 6412 4712 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5994 6440 6000 6452
rect 5031 6412 6000 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 6362 6440 6368 6452
rect 6323 6412 6368 6440
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 15562 6440 15568 6452
rect 6512 6412 15568 6440
rect 6512 6400 6518 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 16022 6440 16028 6452
rect 15983 6412 16028 6440
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16724 6412 17141 6440
rect 16724 6400 16730 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17129 6403 17187 6409
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 19242 6440 19248 6452
rect 17276 6412 19248 6440
rect 17276 6400 17282 6412
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6440 19855 6443
rect 19978 6440 19984 6452
rect 19843 6412 19984 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 22462 6400 22468 6452
rect 22520 6440 22526 6452
rect 27154 6440 27160 6452
rect 22520 6412 27160 6440
rect 22520 6400 22526 6412
rect 27154 6400 27160 6412
rect 27212 6400 27218 6452
rect 27798 6440 27804 6452
rect 27264 6412 27804 6440
rect 8386 6372 8392 6384
rect 5828 6344 8392 6372
rect 5828 6313 5856 6344
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 8938 6372 8944 6384
rect 8899 6344 8944 6372
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 12069 6375 12127 6381
rect 9272 6344 9628 6372
rect 9272 6332 9278 6344
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 6546 6304 6552 6316
rect 6507 6276 6552 6304
rect 5813 6267 5871 6273
rect 4540 6168 4568 6267
rect 5184 6236 5212 6267
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7607 6276 8156 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7282 6236 7288 6248
rect 5184 6208 7288 6236
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 8018 6236 8024 6248
rect 7979 6208 8024 6236
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8128 6236 8156 6276
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 9600 6313 9628 6344
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 12526 6372 12532 6384
rect 12115 6344 12532 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 15933 6375 15991 6381
rect 15933 6372 15945 6375
rect 13596 6344 15945 6372
rect 13596 6332 13602 6344
rect 15933 6341 15945 6344
rect 15979 6341 15991 6375
rect 18684 6375 18742 6381
rect 15933 6335 15991 6341
rect 16592 6344 17816 6372
rect 9585 6307 9643 6313
rect 8260 6276 8305 6304
rect 8260 6264 8266 6276
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 9585 6267 9643 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12980 6307 13038 6313
rect 12980 6273 12992 6307
rect 13026 6304 13038 6307
rect 14550 6304 14556 6316
rect 13026 6276 14412 6304
rect 14511 6276 14556 6304
rect 13026 6273 13038 6276
rect 12980 6267 13038 6273
rect 8938 6236 8944 6248
rect 8128 6208 8944 6236
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9732 6208 9873 6236
rect 9732 6196 9738 6208
rect 9861 6205 9873 6208
rect 9907 6236 9919 6239
rect 9950 6236 9956 6248
rect 9907 6208 9956 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 12710 6236 12716 6248
rect 12671 6208 12716 6236
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 14384 6236 14412 6276
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 14700 6276 14749 6304
rect 14700 6264 14706 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 16592 6304 16620 6344
rect 14976 6276 16620 6304
rect 16669 6307 16727 6313
rect 14976 6264 14982 6276
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 16942 6304 16948 6316
rect 16715 6276 16948 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17788 6313 17816 6344
rect 18684 6341 18696 6375
rect 18730 6372 18742 6375
rect 20254 6372 20260 6384
rect 18730 6344 20260 6372
rect 18730 6341 18742 6344
rect 18684 6335 18742 6341
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 21542 6332 21548 6384
rect 21600 6372 21606 6384
rect 22833 6375 22891 6381
rect 22833 6372 22845 6375
rect 21600 6344 22845 6372
rect 21600 6332 21606 6344
rect 22833 6341 22845 6344
rect 22879 6372 22891 6375
rect 22922 6372 22928 6384
rect 22879 6344 22928 6372
rect 22879 6341 22891 6344
rect 22833 6335 22891 6341
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 26510 6372 26516 6384
rect 26160 6344 26516 6372
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 20441 6307 20499 6313
rect 20441 6273 20453 6307
rect 20487 6304 20499 6307
rect 21560 6304 21588 6332
rect 20487 6276 21588 6304
rect 22097 6307 22155 6313
rect 20487 6273 20499 6276
rect 20441 6267 20499 6273
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 17586 6236 17592 6248
rect 14384 6208 17592 6236
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 18414 6236 18420 6248
rect 18375 6208 18420 6236
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20680 6208 20729 6236
rect 20680 6196 20686 6208
rect 20717 6205 20729 6208
rect 20763 6205 20775 6239
rect 20717 6199 20775 6205
rect 6914 6168 6920 6180
rect 4540 6140 6920 6168
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7377 6171 7435 6177
rect 7377 6137 7389 6171
rect 7423 6168 7435 6171
rect 9030 6168 9036 6180
rect 7423 6140 9036 6168
rect 7423 6137 7435 6140
rect 7377 6131 7435 6137
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 9125 6171 9183 6177
rect 9125 6137 9137 6171
rect 9171 6168 9183 6171
rect 10134 6168 10140 6180
rect 9171 6140 10140 6168
rect 9171 6137 9183 6140
rect 9125 6131 9183 6137
rect 10134 6128 10140 6140
rect 10192 6168 10198 6180
rect 12526 6168 12532 6180
rect 10192 6140 12532 6168
rect 10192 6128 10198 6140
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 18322 6168 18328 6180
rect 16960 6140 18328 6168
rect 5626 6100 5632 6112
rect 5587 6072 5632 6100
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 7524 6072 8401 6100
rect 7524 6060 7530 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 13906 6100 13912 6112
rect 12299 6072 13912 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 16482 6100 16488 6112
rect 14967 6072 16488 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16960 6109 16988 6140
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 20254 6128 20260 6180
rect 20312 6168 20318 6180
rect 21450 6168 21456 6180
rect 20312 6140 21456 6168
rect 20312 6128 20318 6140
rect 21450 6128 21456 6140
rect 21508 6128 21514 6180
rect 22112 6168 22140 6267
rect 22554 6264 22560 6316
rect 22612 6304 22618 6316
rect 22649 6307 22707 6313
rect 22649 6304 22661 6307
rect 22612 6276 22661 6304
rect 22612 6264 22618 6276
rect 22649 6273 22661 6276
rect 22695 6273 22707 6307
rect 22649 6267 22707 6273
rect 23928 6307 23986 6313
rect 23928 6273 23940 6307
rect 23974 6304 23986 6307
rect 24210 6304 24216 6316
rect 23974 6276 24216 6304
rect 23974 6273 23986 6276
rect 23928 6267 23986 6273
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6273 25559 6307
rect 26160 6308 26188 6344
rect 26510 6332 26516 6344
rect 26568 6332 26574 6384
rect 27264 6381 27292 6412
rect 27798 6400 27804 6412
rect 27856 6400 27862 6452
rect 28994 6400 29000 6452
rect 29052 6440 29058 6452
rect 29052 6412 30144 6440
rect 29052 6400 29058 6412
rect 27249 6375 27307 6381
rect 27249 6341 27261 6375
rect 27295 6341 27307 6375
rect 27249 6335 27307 6341
rect 27430 6332 27436 6384
rect 27488 6372 27494 6384
rect 29638 6372 29644 6384
rect 27488 6344 29644 6372
rect 27488 6332 27494 6344
rect 26243 6308 26301 6313
rect 26160 6307 26301 6308
rect 26160 6280 26255 6307
rect 25501 6267 25559 6273
rect 26243 6273 26255 6280
rect 26289 6273 26301 6307
rect 26243 6267 26301 6273
rect 26421 6307 26479 6313
rect 26421 6273 26433 6307
rect 26467 6273 26479 6307
rect 26970 6304 26976 6316
rect 26931 6276 26976 6304
rect 26421 6267 26479 6273
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 25130 6236 25136 6248
rect 25056 6208 25136 6236
rect 23566 6168 23572 6180
rect 22112 6140 23572 6168
rect 23566 6128 23572 6140
rect 23624 6128 23630 6180
rect 25056 6177 25084 6208
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 25516 6236 25544 6267
rect 26436 6236 26464 6267
rect 26970 6264 26976 6276
rect 27028 6264 27034 6316
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 27080 6276 27169 6304
rect 26510 6236 26516 6248
rect 25516 6208 26372 6236
rect 26436 6208 26516 6236
rect 25041 6171 25099 6177
rect 25041 6137 25053 6171
rect 25087 6137 25099 6171
rect 25041 6131 25099 6137
rect 25222 6128 25228 6180
rect 25280 6168 25286 6180
rect 26237 6171 26295 6177
rect 26237 6168 26249 6171
rect 25280 6140 26249 6168
rect 25280 6128 25286 6140
rect 26237 6137 26249 6140
rect 26283 6137 26295 6171
rect 26344 6168 26372 6208
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 26786 6196 26792 6248
rect 26844 6236 26850 6248
rect 27080 6236 27108 6276
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27338 6304 27344 6316
rect 27299 6276 27344 6304
rect 27157 6267 27215 6273
rect 27338 6264 27344 6276
rect 27396 6264 27402 6316
rect 27985 6307 28043 6313
rect 27985 6273 27997 6307
rect 28031 6304 28043 6307
rect 28074 6304 28080 6316
rect 28031 6276 28080 6304
rect 28031 6273 28043 6276
rect 27985 6267 28043 6273
rect 28074 6264 28080 6276
rect 28132 6264 28138 6316
rect 28169 6307 28227 6313
rect 28169 6273 28181 6307
rect 28215 6273 28227 6307
rect 28169 6267 28227 6273
rect 28184 6236 28212 6267
rect 28258 6264 28264 6316
rect 28316 6304 28322 6316
rect 28399 6307 28457 6313
rect 28316 6276 28361 6304
rect 28316 6264 28322 6276
rect 28399 6273 28411 6307
rect 28445 6304 28457 6307
rect 28534 6304 28540 6316
rect 28445 6276 28540 6304
rect 28445 6273 28457 6276
rect 28399 6267 28457 6273
rect 28534 6264 28540 6276
rect 28592 6264 28598 6316
rect 29104 6313 29132 6344
rect 29638 6332 29644 6344
rect 29696 6332 29702 6384
rect 30116 6372 30144 6412
rect 30190 6400 30196 6452
rect 30248 6440 30254 6452
rect 30469 6443 30527 6449
rect 30469 6440 30481 6443
rect 30248 6412 30481 6440
rect 30248 6400 30254 6412
rect 30469 6409 30481 6412
rect 30515 6409 30527 6443
rect 34701 6443 34759 6449
rect 30469 6403 30527 6409
rect 31726 6412 34376 6440
rect 30282 6372 30288 6384
rect 30116 6344 30288 6372
rect 30282 6332 30288 6344
rect 30340 6372 30346 6384
rect 30340 6344 31156 6372
rect 30340 6332 30346 6344
rect 29362 6313 29368 6316
rect 29089 6307 29147 6313
rect 29089 6273 29101 6307
rect 29135 6273 29147 6307
rect 29356 6304 29368 6313
rect 29323 6276 29368 6304
rect 29089 6267 29147 6273
rect 29356 6267 29368 6276
rect 29362 6264 29368 6267
rect 29420 6264 29426 6316
rect 30374 6264 30380 6316
rect 30432 6304 30438 6316
rect 31128 6313 31156 6344
rect 30929 6307 30987 6313
rect 30929 6304 30941 6307
rect 30432 6276 30941 6304
rect 30432 6264 30438 6276
rect 30929 6273 30941 6276
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6273 31171 6307
rect 31113 6267 31171 6273
rect 26844 6208 28672 6236
rect 26844 6196 26850 6208
rect 26694 6168 26700 6180
rect 26344 6140 26700 6168
rect 26237 6131 26295 6137
rect 26694 6128 26700 6140
rect 26752 6128 26758 6180
rect 28442 6168 28448 6180
rect 27356 6140 28448 6168
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6069 17003 6103
rect 16945 6063 17003 6069
rect 17494 6060 17500 6112
rect 17552 6100 17558 6112
rect 17589 6103 17647 6109
rect 17589 6100 17601 6103
rect 17552 6072 17601 6100
rect 17552 6060 17558 6072
rect 17589 6069 17601 6072
rect 17635 6069 17647 6103
rect 17589 6063 17647 6069
rect 21913 6103 21971 6109
rect 21913 6069 21925 6103
rect 21959 6100 21971 6103
rect 22646 6100 22652 6112
rect 21959 6072 22652 6100
rect 21959 6069 21971 6072
rect 21913 6063 21971 6069
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 23382 6060 23388 6112
rect 23440 6100 23446 6112
rect 25685 6103 25743 6109
rect 25685 6100 25697 6103
rect 23440 6072 25697 6100
rect 23440 6060 23446 6072
rect 25685 6069 25697 6072
rect 25731 6069 25743 6103
rect 25685 6063 25743 6069
rect 25958 6060 25964 6112
rect 26016 6100 26022 6112
rect 27356 6100 27384 6140
rect 28442 6128 28448 6140
rect 28500 6128 28506 6180
rect 26016 6072 27384 6100
rect 26016 6060 26022 6072
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 27525 6103 27583 6109
rect 27525 6100 27537 6103
rect 27488 6072 27537 6100
rect 27488 6060 27494 6072
rect 27525 6069 27537 6072
rect 27571 6069 27583 6103
rect 27525 6063 27583 6069
rect 28350 6060 28356 6112
rect 28408 6100 28414 6112
rect 28537 6103 28595 6109
rect 28537 6100 28549 6103
rect 28408 6072 28549 6100
rect 28408 6060 28414 6072
rect 28537 6069 28549 6072
rect 28583 6069 28595 6103
rect 28644 6100 28672 6208
rect 31726 6168 31754 6412
rect 32030 6332 32036 6384
rect 32088 6372 32094 6384
rect 32309 6375 32367 6381
rect 32309 6372 32321 6375
rect 32088 6344 32321 6372
rect 32088 6332 32094 6344
rect 32309 6341 32321 6344
rect 32355 6372 32367 6375
rect 33042 6372 33048 6384
rect 32355 6344 33048 6372
rect 32355 6341 32367 6344
rect 32309 6335 32367 6341
rect 33042 6332 33048 6344
rect 33100 6332 33106 6384
rect 34348 6381 34376 6412
rect 34701 6409 34713 6443
rect 34747 6440 34759 6443
rect 34790 6440 34796 6452
rect 34747 6412 34796 6440
rect 34747 6409 34759 6412
rect 34701 6403 34759 6409
rect 34790 6400 34796 6412
rect 34848 6400 34854 6452
rect 35158 6400 35164 6452
rect 35216 6440 35222 6452
rect 35618 6440 35624 6452
rect 35216 6412 35624 6440
rect 35216 6400 35222 6412
rect 35618 6400 35624 6412
rect 35676 6400 35682 6452
rect 35713 6443 35771 6449
rect 35713 6409 35725 6443
rect 35759 6409 35771 6443
rect 35713 6403 35771 6409
rect 34333 6375 34391 6381
rect 34333 6341 34345 6375
rect 34379 6372 34391 6375
rect 35066 6372 35072 6384
rect 34379 6344 35072 6372
rect 34379 6341 34391 6344
rect 34333 6335 34391 6341
rect 35066 6332 35072 6344
rect 35124 6372 35130 6384
rect 35345 6375 35403 6381
rect 35345 6372 35357 6375
rect 35124 6344 35357 6372
rect 35124 6332 35130 6344
rect 35345 6341 35357 6344
rect 35391 6341 35403 6375
rect 35345 6335 35403 6341
rect 35437 6375 35495 6381
rect 35437 6341 35449 6375
rect 35483 6372 35495 6375
rect 35483 6344 35664 6372
rect 35483 6341 35495 6344
rect 35437 6335 35495 6341
rect 35636 6316 35664 6344
rect 35728 6316 35756 6403
rect 35802 6400 35808 6452
rect 35860 6440 35866 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 35860 6412 36553 6440
rect 35860 6400 35866 6412
rect 36541 6409 36553 6412
rect 36587 6409 36599 6443
rect 36541 6403 36599 6409
rect 36173 6375 36231 6381
rect 36173 6341 36185 6375
rect 36219 6372 36231 6375
rect 36262 6372 36268 6384
rect 36219 6344 36268 6372
rect 36219 6341 36231 6344
rect 36173 6335 36231 6341
rect 36262 6332 36268 6344
rect 36320 6332 36326 6384
rect 32125 6307 32183 6313
rect 32125 6273 32137 6307
rect 32171 6304 32183 6307
rect 32674 6304 32680 6316
rect 32171 6276 32680 6304
rect 32171 6273 32183 6276
rect 32125 6267 32183 6273
rect 32674 6264 32680 6276
rect 32732 6264 32738 6316
rect 33134 6304 33140 6316
rect 33095 6276 33140 6304
rect 33134 6264 33140 6276
rect 33192 6264 33198 6316
rect 33686 6264 33692 6316
rect 33744 6304 33750 6316
rect 34149 6307 34207 6313
rect 34149 6304 34161 6307
rect 33744 6276 34161 6304
rect 33744 6264 33750 6276
rect 34149 6273 34161 6276
rect 34195 6273 34207 6307
rect 34149 6267 34207 6273
rect 34238 6264 34244 6316
rect 34296 6304 34302 6316
rect 34425 6307 34483 6313
rect 34425 6304 34437 6307
rect 34296 6276 34437 6304
rect 34296 6264 34302 6276
rect 34425 6273 34437 6276
rect 34471 6273 34483 6307
rect 34425 6267 34483 6273
rect 34517 6307 34575 6313
rect 34517 6273 34529 6307
rect 34563 6273 34575 6307
rect 35158 6304 35164 6316
rect 35119 6276 35164 6304
rect 34517 6267 34575 6273
rect 32493 6239 32551 6245
rect 32493 6205 32505 6239
rect 32539 6236 32551 6239
rect 34532 6236 34560 6267
rect 35158 6264 35164 6276
rect 35216 6264 35222 6316
rect 35529 6307 35587 6313
rect 35529 6304 35541 6307
rect 35360 6276 35541 6304
rect 35360 6248 35388 6276
rect 35529 6273 35541 6276
rect 35575 6273 35587 6307
rect 35529 6267 35587 6273
rect 35618 6264 35624 6316
rect 35676 6264 35682 6316
rect 35710 6264 35716 6316
rect 35768 6264 35774 6316
rect 36357 6307 36415 6313
rect 36357 6273 36369 6307
rect 36403 6273 36415 6307
rect 36357 6267 36415 6273
rect 35342 6236 35348 6248
rect 32539 6208 34376 6236
rect 34532 6208 35348 6236
rect 32539 6205 32551 6208
rect 32493 6199 32551 6205
rect 30024 6140 31754 6168
rect 30024 6100 30052 6140
rect 31938 6128 31944 6180
rect 31996 6168 32002 6180
rect 32953 6171 33011 6177
rect 32953 6168 32965 6171
rect 31996 6140 32965 6168
rect 31996 6128 32002 6140
rect 32953 6137 32965 6140
rect 32999 6137 33011 6171
rect 34348 6168 34376 6208
rect 35342 6196 35348 6208
rect 35400 6196 35406 6248
rect 35452 6208 35848 6236
rect 35452 6168 35480 6208
rect 34348 6140 35480 6168
rect 35820 6168 35848 6208
rect 35986 6196 35992 6248
rect 36044 6236 36050 6248
rect 36372 6236 36400 6267
rect 36044 6208 36400 6236
rect 36044 6196 36050 6208
rect 36170 6168 36176 6180
rect 35820 6140 36176 6168
rect 32953 6131 33011 6137
rect 36170 6128 36176 6140
rect 36228 6128 36234 6180
rect 28644 6072 30052 6100
rect 30929 6103 30987 6109
rect 28537 6063 28595 6069
rect 30929 6069 30941 6103
rect 30975 6100 30987 6103
rect 37458 6100 37464 6112
rect 30975 6072 37464 6100
rect 30975 6069 30987 6072
rect 30929 6063 30987 6069
rect 37458 6060 37464 6072
rect 37516 6060 37522 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 5074 5896 5080 5908
rect 5035 5868 5080 5896
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 5684 5868 11744 5896
rect 5684 5856 5690 5868
rect 5721 5831 5779 5837
rect 5721 5797 5733 5831
rect 5767 5828 5779 5831
rect 6454 5828 6460 5840
rect 5767 5800 6460 5828
rect 5767 5797 5779 5800
rect 5721 5791 5779 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7558 5828 7564 5840
rect 6972 5800 7564 5828
rect 6972 5788 6978 5800
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 11716 5828 11744 5868
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 11940 5868 13001 5896
rect 11940 5856 11946 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 12989 5859 13047 5865
rect 13449 5899 13507 5905
rect 13449 5865 13461 5899
rect 13495 5896 13507 5899
rect 13722 5896 13728 5908
rect 13495 5868 13728 5896
rect 13495 5865 13507 5868
rect 13449 5859 13507 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14918 5896 14924 5908
rect 13872 5868 14924 5896
rect 13872 5856 13878 5868
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 17586 5896 17592 5908
rect 15896 5868 17448 5896
rect 17547 5868 17592 5896
rect 15896 5856 15902 5868
rect 11716 5800 13584 5828
rect 8297 5763 8355 5769
rect 8297 5760 8309 5763
rect 6564 5732 8309 5760
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5718 5692 5724 5704
rect 5307 5664 5724 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 6564 5701 6592 5732
rect 8297 5729 8309 5732
rect 8343 5729 8355 5763
rect 8297 5723 8355 5729
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 7466 5692 7472 5704
rect 7427 5664 7472 5692
rect 6549 5655 6607 5661
rect 5920 5624 5948 5655
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8754 5692 8760 5704
rect 8159 5664 8760 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 8987 5664 10793 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 10781 5661 10793 5664
rect 10827 5692 10839 5695
rect 12158 5692 12164 5704
rect 10827 5664 12164 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 6730 5624 6736 5636
rect 5920 5596 6736 5624
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 6822 5584 6828 5636
rect 6880 5624 6886 5636
rect 8956 5624 8984 5655
rect 12158 5652 12164 5664
rect 12216 5692 12222 5704
rect 12710 5692 12716 5704
rect 12216 5664 12716 5692
rect 12216 5652 12222 5664
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 13170 5692 13176 5704
rect 13131 5664 13176 5692
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13556 5701 13584 5800
rect 13906 5788 13912 5840
rect 13964 5828 13970 5840
rect 16025 5831 16083 5837
rect 13964 5800 15700 5828
rect 13964 5788 13970 5800
rect 14734 5760 14740 5772
rect 14695 5732 14740 5760
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 15672 5760 15700 5800
rect 16025 5797 16037 5831
rect 16071 5828 16083 5831
rect 16298 5828 16304 5840
rect 16071 5800 16304 5828
rect 16071 5797 16083 5800
rect 16025 5791 16083 5797
rect 16298 5788 16304 5800
rect 16356 5788 16362 5840
rect 16942 5828 16948 5840
rect 16903 5800 16948 5828
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17037 5831 17095 5837
rect 17037 5797 17049 5831
rect 17083 5828 17095 5831
rect 17310 5828 17316 5840
rect 17083 5800 17316 5828
rect 17083 5797 17095 5800
rect 17037 5791 17095 5797
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 17420 5828 17448 5868
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 20530 5896 20536 5908
rect 17696 5868 20536 5896
rect 17696 5828 17724 5868
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 21910 5896 21916 5908
rect 21871 5868 21916 5896
rect 21910 5856 21916 5868
rect 21968 5856 21974 5908
rect 26050 5896 26056 5908
rect 22066 5868 25636 5896
rect 26011 5868 26056 5896
rect 17420 5800 17724 5828
rect 18414 5788 18420 5840
rect 18472 5788 18478 5840
rect 19334 5788 19340 5840
rect 19392 5828 19398 5840
rect 19429 5831 19487 5837
rect 19429 5828 19441 5831
rect 19392 5800 19441 5828
rect 19392 5788 19398 5800
rect 19429 5797 19441 5800
rect 19475 5797 19487 5831
rect 22066 5828 22094 5868
rect 19429 5791 19487 5797
rect 21560 5800 22094 5828
rect 25608 5828 25636 5868
rect 26050 5856 26056 5868
rect 26108 5856 26114 5908
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 27893 5899 27951 5905
rect 27893 5896 27905 5899
rect 27856 5868 27905 5896
rect 27856 5856 27862 5868
rect 27893 5865 27905 5868
rect 27939 5865 27951 5899
rect 27893 5859 27951 5865
rect 28000 5868 31800 5896
rect 25958 5828 25964 5840
rect 25608 5800 25964 5828
rect 18432 5760 18460 5788
rect 20530 5760 20536 5772
rect 15672 5732 17816 5760
rect 18432 5732 20536 5760
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 6880 5596 8984 5624
rect 6880 5584 6886 5596
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9186 5627 9244 5633
rect 9186 5624 9198 5627
rect 9088 5596 9198 5624
rect 9088 5584 9094 5596
rect 9186 5593 9198 5596
rect 9232 5593 9244 5627
rect 9186 5587 9244 5593
rect 11048 5627 11106 5633
rect 11048 5593 11060 5627
rect 11094 5624 11106 5627
rect 12342 5624 12348 5636
rect 11094 5596 12348 5624
rect 11094 5593 11106 5596
rect 11048 5587 11106 5593
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 13280 5624 13308 5655
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14148 5664 14657 5692
rect 14148 5652 14154 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14884 5664 14933 5692
rect 14884 5652 14890 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 14921 5655 14979 5661
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 17310 5692 17316 5704
rect 16071 5664 17316 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 14108 5624 14136 5652
rect 13280 5596 14136 5624
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 15010 5624 15016 5636
rect 14240 5596 15016 5624
rect 14240 5584 14246 5596
rect 15010 5584 15016 5596
rect 15068 5624 15074 5636
rect 16040 5624 16068 5655
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17788 5701 17816 5732
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18288 5664 18429 5692
rect 18288 5652 18294 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18966 5652 18972 5704
rect 19024 5692 19030 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19024 5664 19257 5692
rect 19024 5652 19030 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 19245 5655 19303 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5692 20131 5695
rect 20162 5692 20168 5704
rect 20119 5664 20168 5692
rect 20119 5661 20131 5664
rect 20073 5655 20131 5661
rect 15068 5596 16068 5624
rect 16577 5627 16635 5633
rect 15068 5584 15074 5596
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 18322 5624 18328 5636
rect 16623 5596 18328 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 18322 5584 18328 5596
rect 18380 5584 18386 5636
rect 19812 5624 19840 5655
rect 20162 5652 20168 5664
rect 20220 5692 20226 5704
rect 21560 5692 21588 5800
rect 25958 5788 25964 5800
rect 26016 5788 26022 5840
rect 27614 5788 27620 5840
rect 27672 5828 27678 5840
rect 28000 5828 28028 5868
rect 27672 5800 28028 5828
rect 31772 5828 31800 5868
rect 34238 5856 34244 5908
rect 34296 5896 34302 5908
rect 36081 5899 36139 5905
rect 36081 5896 36093 5899
rect 34296 5868 36093 5896
rect 34296 5856 34302 5868
rect 36081 5865 36093 5868
rect 36127 5865 36139 5899
rect 36081 5859 36139 5865
rect 36170 5856 36176 5908
rect 36228 5896 36234 5908
rect 37185 5899 37243 5905
rect 37185 5896 37197 5899
rect 36228 5868 37197 5896
rect 36228 5856 36234 5868
rect 37185 5865 37197 5868
rect 37231 5865 37243 5899
rect 37185 5859 37243 5865
rect 33505 5831 33563 5837
rect 33505 5828 33517 5831
rect 31772 5800 33517 5828
rect 27672 5788 27678 5800
rect 33505 5797 33517 5800
rect 33551 5797 33563 5831
rect 33505 5791 33563 5797
rect 36541 5831 36599 5837
rect 36541 5797 36553 5831
rect 36587 5828 36599 5831
rect 37826 5828 37832 5840
rect 36587 5800 37832 5828
rect 36587 5797 36599 5800
rect 36541 5791 36599 5797
rect 37826 5788 37832 5800
rect 37884 5788 37890 5840
rect 22554 5760 22560 5772
rect 22515 5732 22560 5760
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 22833 5763 22891 5769
rect 22833 5729 22845 5763
rect 22879 5760 22891 5763
rect 23014 5760 23020 5772
rect 22879 5732 23020 5760
rect 22879 5729 22891 5732
rect 22833 5723 22891 5729
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 29822 5760 29828 5772
rect 27632 5732 28994 5760
rect 29783 5732 29828 5760
rect 20220 5664 21588 5692
rect 20220 5652 20226 5664
rect 23658 5652 23664 5704
rect 23716 5692 23722 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 23716 5664 24685 5692
rect 23716 5652 23722 5664
rect 24673 5661 24685 5664
rect 24719 5692 24731 5695
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 24719 5664 26525 5692
rect 24719 5661 24731 5664
rect 24673 5655 24731 5661
rect 26513 5661 26525 5664
rect 26559 5692 26571 5695
rect 27246 5692 27252 5704
rect 26559 5664 27252 5692
rect 26559 5661 26571 5664
rect 26513 5655 26571 5661
rect 27246 5652 27252 5664
rect 27304 5652 27310 5704
rect 20622 5624 20628 5636
rect 19812 5596 20628 5624
rect 20622 5584 20628 5596
rect 20680 5584 20686 5636
rect 20800 5627 20858 5633
rect 20800 5593 20812 5627
rect 20846 5624 20858 5627
rect 20898 5624 20904 5636
rect 20846 5596 20904 5624
rect 20846 5593 20858 5596
rect 20800 5587 20858 5593
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 24940 5627 24998 5633
rect 24940 5593 24952 5627
rect 24986 5624 24998 5627
rect 25682 5624 25688 5636
rect 24986 5596 25688 5624
rect 24986 5593 24998 5596
rect 24940 5587 24998 5593
rect 25682 5584 25688 5596
rect 25740 5584 25746 5636
rect 26234 5584 26240 5636
rect 26292 5624 26298 5636
rect 26758 5627 26816 5633
rect 26758 5624 26770 5627
rect 26292 5596 26770 5624
rect 26292 5584 26298 5596
rect 26758 5593 26770 5596
rect 26804 5593 26816 5627
rect 26758 5587 26816 5593
rect 26878 5584 26884 5636
rect 26936 5624 26942 5636
rect 27632 5624 27660 5732
rect 28074 5652 28080 5704
rect 28132 5692 28138 5704
rect 28534 5692 28540 5704
rect 28132 5664 28540 5692
rect 28132 5652 28138 5664
rect 28534 5652 28540 5664
rect 28592 5652 28598 5704
rect 28966 5692 28994 5732
rect 29822 5720 29828 5732
rect 29880 5720 29886 5772
rect 32122 5760 32128 5772
rect 30852 5732 32128 5760
rect 30852 5692 30880 5732
rect 32122 5720 32128 5732
rect 32180 5720 32186 5772
rect 32582 5720 32588 5772
rect 32640 5760 32646 5772
rect 34698 5760 34704 5772
rect 32640 5732 34560 5760
rect 34659 5732 34704 5760
rect 32640 5720 32646 5732
rect 28966 5664 30880 5692
rect 31018 5652 31024 5704
rect 31076 5692 31082 5704
rect 31665 5695 31723 5701
rect 31665 5692 31677 5695
rect 31076 5664 31677 5692
rect 31076 5652 31082 5664
rect 31665 5661 31677 5664
rect 31711 5661 31723 5695
rect 31665 5655 31723 5661
rect 31754 5652 31760 5704
rect 31812 5692 31818 5704
rect 31849 5695 31907 5701
rect 31849 5692 31861 5695
rect 31812 5664 31861 5692
rect 31812 5652 31818 5664
rect 31849 5661 31861 5664
rect 31895 5661 31907 5695
rect 33410 5692 33416 5704
rect 31849 5655 31907 5661
rect 32508 5664 33416 5692
rect 28994 5624 29000 5636
rect 26936 5596 27660 5624
rect 27688 5596 29000 5624
rect 26936 5584 26942 5596
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6454 5556 6460 5568
rect 6411 5528 6460 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 7156 5528 7297 5556
rect 7156 5516 7162 5528
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7285 5519 7343 5525
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8294 5556 8300 5568
rect 8076 5528 8300 5556
rect 8076 5516 8082 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 10284 5528 10333 5556
rect 10284 5516 10290 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 10321 5519 10379 5525
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11848 5528 12173 5556
rect 11848 5516 11854 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 16298 5556 16304 5568
rect 15160 5528 16304 5556
rect 15160 5516 15166 5528
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 18598 5556 18604 5568
rect 18559 5528 18604 5556
rect 18598 5516 18604 5528
rect 18656 5556 18662 5568
rect 23106 5556 23112 5568
rect 18656 5528 23112 5556
rect 18656 5516 18662 5528
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 26510 5516 26516 5568
rect 26568 5556 26574 5568
rect 27688 5556 27716 5596
rect 28994 5584 29000 5596
rect 29052 5584 29058 5636
rect 30092 5627 30150 5633
rect 30092 5593 30104 5627
rect 30138 5624 30150 5627
rect 32508 5624 32536 5664
rect 33410 5652 33416 5664
rect 33468 5652 33474 5704
rect 33686 5692 33692 5704
rect 33647 5664 33692 5692
rect 33686 5652 33692 5664
rect 33744 5652 33750 5704
rect 34532 5692 34560 5732
rect 34698 5720 34704 5732
rect 34756 5720 34762 5772
rect 36188 5732 38056 5760
rect 34606 5692 34612 5704
rect 34532 5664 34612 5692
rect 34606 5652 34612 5664
rect 34664 5652 34670 5704
rect 36188 5692 36216 5732
rect 34900 5664 36216 5692
rect 32674 5624 32680 5636
rect 30138 5596 32536 5624
rect 32587 5596 32680 5624
rect 30138 5593 30150 5596
rect 30092 5587 30150 5593
rect 32674 5584 32680 5596
rect 32732 5584 32738 5636
rect 32858 5624 32864 5636
rect 32819 5596 32864 5624
rect 32858 5584 32864 5596
rect 32916 5584 32922 5636
rect 33045 5627 33103 5633
rect 33045 5593 33057 5627
rect 33091 5624 33103 5627
rect 34900 5624 34928 5664
rect 36722 5652 36728 5704
rect 36780 5652 36786 5704
rect 38028 5701 38056 5732
rect 37369 5695 37427 5701
rect 37369 5692 37381 5695
rect 36832 5664 37381 5692
rect 36725 5637 36737 5652
rect 36771 5637 36783 5652
rect 33091 5596 34928 5624
rect 34968 5627 35026 5633
rect 33091 5593 33103 5596
rect 33045 5587 33103 5593
rect 34968 5593 34980 5627
rect 35014 5624 35026 5627
rect 36078 5624 36084 5636
rect 35014 5596 36084 5624
rect 35014 5593 35026 5596
rect 34968 5587 35026 5593
rect 36078 5584 36084 5596
rect 36136 5584 36142 5636
rect 36725 5631 36783 5637
rect 26568 5528 27716 5556
rect 26568 5516 26574 5528
rect 27798 5516 27804 5568
rect 27856 5556 27862 5568
rect 28353 5559 28411 5565
rect 28353 5556 28365 5559
rect 27856 5528 28365 5556
rect 27856 5516 27862 5528
rect 28353 5525 28365 5528
rect 28399 5525 28411 5559
rect 28353 5519 28411 5525
rect 30834 5516 30840 5568
rect 30892 5556 30898 5568
rect 31205 5559 31263 5565
rect 31205 5556 31217 5559
rect 30892 5528 31217 5556
rect 30892 5516 30898 5528
rect 31205 5525 31217 5528
rect 31251 5525 31263 5559
rect 31205 5519 31263 5525
rect 31757 5559 31815 5565
rect 31757 5525 31769 5559
rect 31803 5556 31815 5559
rect 32582 5556 32588 5568
rect 31803 5528 32588 5556
rect 31803 5525 31815 5528
rect 31757 5519 31815 5525
rect 32582 5516 32588 5528
rect 32640 5516 32646 5568
rect 32692 5556 32720 5584
rect 33870 5556 33876 5568
rect 32692 5528 33876 5556
rect 33870 5516 33876 5528
rect 33928 5516 33934 5568
rect 34238 5516 34244 5568
rect 34296 5556 34302 5568
rect 36832 5556 36860 5664
rect 37369 5661 37381 5664
rect 37415 5661 37427 5695
rect 37369 5655 37427 5661
rect 38013 5695 38071 5701
rect 38013 5661 38025 5695
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 34296 5528 36860 5556
rect 34296 5516 34302 5528
rect 36906 5516 36912 5568
rect 36964 5556 36970 5568
rect 37829 5559 37887 5565
rect 37829 5556 37841 5559
rect 36964 5528 37841 5556
rect 36964 5516 36970 5528
rect 37829 5525 37841 5528
rect 37875 5525 37887 5559
rect 37829 5519 37887 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 5442 5352 5448 5364
rect 4203 5324 5448 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 8754 5352 8760 5364
rect 5684 5324 8524 5352
rect 8715 5324 8760 5352
rect 5684 5312 5690 5324
rect 5994 5284 6000 5296
rect 4356 5256 6000 5284
rect 4356 5225 4384 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 6822 5284 6828 5296
rect 6380 5256 6828 5284
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 5902 5216 5908 5228
rect 5859 5188 5908 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 5184 5148 5212 5179
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6380 5225 6408 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 8018 5284 8024 5296
rect 6972 5256 8024 5284
rect 6972 5244 6978 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8496 5293 8524 5324
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9048 5324 9628 5352
rect 8481 5287 8539 5293
rect 8481 5253 8493 5287
rect 8527 5253 8539 5287
rect 9048 5284 9076 5324
rect 8481 5247 8539 5253
rect 8588 5256 9076 5284
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6621 5219 6679 5225
rect 6621 5216 6633 5219
rect 6512 5188 6633 5216
rect 6512 5176 6518 5188
rect 6621 5185 6633 5188
rect 6667 5185 6679 5219
rect 6621 5179 6679 5185
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8588 5225 8616 5256
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9401 5287 9459 5293
rect 9401 5284 9413 5287
rect 9180 5256 9413 5284
rect 9180 5244 9186 5256
rect 9401 5253 9413 5256
rect 9447 5253 9459 5287
rect 9401 5247 9459 5253
rect 9600 5284 9628 5324
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 9732 5324 10456 5352
rect 9732 5312 9738 5324
rect 10042 5284 10048 5296
rect 9600 5256 10048 5284
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7892 5188 8217 5216
rect 7892 5176 7898 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 6086 5148 6092 5160
rect 4755 5120 6092 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 8404 5148 8432 5179
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 9600 5225 9628 5256
rect 10042 5244 10048 5256
rect 10100 5284 10106 5296
rect 10428 5293 10456 5324
rect 10594 5312 10600 5364
rect 10652 5312 10658 5364
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 14550 5352 14556 5364
rect 13403 5324 14556 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 14976 5324 15761 5352
rect 14976 5312 14982 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 15749 5315 15807 5321
rect 18141 5355 18199 5361
rect 18141 5321 18153 5355
rect 18187 5352 18199 5355
rect 18322 5352 18328 5364
rect 18187 5324 18328 5352
rect 18187 5321 18199 5324
rect 18141 5315 18199 5321
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 22462 5352 22468 5364
rect 20588 5324 22468 5352
rect 20588 5312 20594 5324
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 23014 5352 23020 5364
rect 22572 5324 23020 5352
rect 10413 5287 10471 5293
rect 10100 5256 10364 5284
rect 10100 5244 10106 5256
rect 9237 5219 9295 5225
rect 9237 5216 9249 5219
rect 8720 5188 9249 5216
rect 8720 5176 8726 5188
rect 9237 5185 9249 5188
rect 9283 5185 9295 5219
rect 9237 5179 9295 5185
rect 9489 5219 9547 5225
rect 9489 5212 9501 5219
rect 9535 5212 9547 5219
rect 9585 5219 9643 5225
rect 9489 5179 9496 5212
rect 9490 5160 9496 5179
rect 9548 5160 9554 5212
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 10226 5216 10232 5228
rect 10187 5188 10232 5216
rect 9585 5179 9643 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10336 5216 10364 5256
rect 10413 5253 10425 5287
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 10505 5287 10563 5293
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 10612 5284 10640 5312
rect 13170 5284 13176 5296
rect 10551 5256 10640 5284
rect 11716 5256 13176 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 11716 5225 11744 5256
rect 13170 5244 13176 5256
rect 13228 5284 13234 5296
rect 15194 5284 15200 5296
rect 13228 5256 13584 5284
rect 13228 5244 13234 5256
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10336 5188 10609 5216
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12066 5216 12072 5228
rect 11848 5188 11893 5216
rect 12027 5188 12072 5216
rect 11848 5176 11854 5188
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12406 5188 12541 5216
rect 9122 5148 9128 5160
rect 8404 5120 9128 5148
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 12406 5148 12434 5188
rect 12529 5185 12541 5188
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 12802 5216 12808 5228
rect 12759 5188 12808 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13556 5225 13584 5256
rect 14384 5256 15200 5284
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 13814 5216 13820 5228
rect 13679 5188 13820 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14384 5225 14412 5256
rect 15194 5244 15200 5256
rect 15252 5284 15258 5296
rect 16022 5284 16028 5296
rect 15252 5256 16028 5284
rect 15252 5244 15258 5256
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 18414 5284 18420 5296
rect 16776 5256 18420 5284
rect 14369 5219 14427 5225
rect 13964 5188 14009 5216
rect 13964 5176 13970 5188
rect 14369 5185 14381 5219
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 14636 5219 14694 5225
rect 14636 5185 14648 5219
rect 14682 5216 14694 5219
rect 15930 5216 15936 5228
rect 14682 5188 15936 5216
rect 14682 5185 14694 5188
rect 14636 5179 14694 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16040 5216 16068 5244
rect 16776 5225 16804 5256
rect 18414 5244 18420 5256
rect 18472 5244 18478 5296
rect 21913 5287 21971 5293
rect 19076 5256 20386 5284
rect 19076 5228 19104 5256
rect 17034 5225 17040 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16040 5188 16773 5216
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 17028 5179 17040 5225
rect 17092 5216 17098 5228
rect 18782 5216 18788 5228
rect 17092 5188 17128 5216
rect 18743 5188 18788 5216
rect 17034 5176 17040 5179
rect 17092 5176 17098 5188
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5216 19027 5219
rect 19058 5216 19064 5228
rect 19015 5188 19064 5216
rect 19015 5185 19027 5188
rect 18969 5179 19027 5185
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 20165 5219 20223 5225
rect 19659 5188 20116 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 10836 5120 12434 5148
rect 20088 5148 20116 5188
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 20254 5216 20260 5228
rect 20211 5188 20260 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20358 5225 20386 5256
rect 21913 5253 21925 5287
rect 21959 5284 21971 5287
rect 22572 5284 22600 5324
rect 23014 5312 23020 5324
rect 23072 5312 23078 5364
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 25041 5355 25099 5361
rect 25041 5352 25053 5355
rect 23164 5324 25053 5352
rect 23164 5312 23170 5324
rect 25041 5321 25053 5324
rect 25087 5321 25099 5355
rect 26418 5352 26424 5364
rect 26379 5324 26424 5352
rect 25041 5315 25099 5321
rect 26418 5312 26424 5324
rect 26476 5312 26482 5364
rect 27430 5352 27436 5364
rect 27080 5324 27436 5352
rect 21959 5256 22600 5284
rect 21959 5253 21971 5256
rect 21913 5247 21971 5253
rect 22646 5244 22652 5296
rect 22704 5284 22710 5296
rect 26237 5287 26295 5293
rect 22704 5256 24900 5284
rect 22704 5244 22710 5256
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5185 20407 5219
rect 20349 5179 20407 5185
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 20898 5148 20904 5160
rect 20088 5120 20904 5148
rect 10836 5108 10842 5120
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 21008 5148 21036 5179
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22152 5188 22197 5216
rect 22152 5176 22158 5188
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 23290 5216 23296 5228
rect 22336 5188 22381 5216
rect 23251 5188 23296 5216
rect 22336 5176 22342 5188
rect 23290 5176 23296 5188
rect 23348 5176 23354 5228
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5216 23443 5219
rect 23474 5216 23480 5228
rect 23431 5188 23480 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5216 23719 5219
rect 23842 5216 23848 5228
rect 23707 5188 23848 5216
rect 23707 5185 23719 5188
rect 23661 5179 23719 5185
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24872 5225 24900 5256
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 27080 5284 27108 5324
rect 27430 5312 27436 5324
rect 27488 5312 27494 5364
rect 28258 5312 28264 5364
rect 28316 5352 28322 5364
rect 28629 5355 28687 5361
rect 28629 5352 28641 5355
rect 28316 5324 28641 5352
rect 28316 5312 28322 5324
rect 28629 5321 28641 5324
rect 28675 5321 28687 5355
rect 33226 5352 33232 5364
rect 28629 5315 28687 5321
rect 28736 5324 33232 5352
rect 27614 5284 27620 5296
rect 26283 5256 27108 5284
rect 27264 5256 27620 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 27264 5228 27292 5256
rect 27614 5244 27620 5256
rect 27672 5244 27678 5296
rect 27706 5244 27712 5296
rect 27764 5284 27770 5296
rect 28736 5284 28764 5324
rect 33226 5312 33232 5324
rect 33284 5312 33290 5364
rect 34238 5352 34244 5364
rect 34199 5324 34244 5352
rect 34238 5312 34244 5324
rect 34296 5312 34302 5364
rect 35618 5312 35624 5364
rect 35676 5352 35682 5364
rect 36081 5355 36139 5361
rect 36081 5352 36093 5355
rect 35676 5324 36093 5352
rect 35676 5312 35682 5324
rect 36081 5321 36093 5324
rect 36127 5321 36139 5355
rect 36081 5315 36139 5321
rect 31294 5284 31300 5296
rect 27764 5256 28764 5284
rect 30392 5256 31300 5284
rect 27764 5244 27770 5256
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 24176 5188 24225 5216
rect 24176 5176 24182 5188
rect 24213 5185 24225 5188
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24857 5219 24915 5225
rect 24857 5185 24869 5219
rect 24903 5185 24915 5219
rect 24857 5179 24915 5185
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5216 26111 5219
rect 27246 5216 27252 5228
rect 26099 5188 27108 5216
rect 27207 5188 27252 5216
rect 26099 5185 26111 5188
rect 26053 5179 26111 5185
rect 22186 5148 22192 5160
rect 21008 5120 22192 5148
rect 22186 5108 22192 5120
rect 22244 5108 22250 5160
rect 26418 5108 26424 5160
rect 26476 5148 26482 5160
rect 26878 5148 26884 5160
rect 26476 5120 26884 5148
rect 26476 5108 26482 5120
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 6362 5080 6368 5092
rect 6012 5052 6368 5080
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3568 4984 3801 5012
rect 3568 4972 3574 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 3789 4975 3847 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 6012 5012 6040 5052
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 10410 5080 10416 5092
rect 7300 5052 10416 5080
rect 5675 4984 6040 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 7300 5012 7328 5052
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 10870 5040 10876 5092
rect 10928 5080 10934 5092
rect 11977 5083 12035 5089
rect 11977 5080 11989 5083
rect 10928 5052 11989 5080
rect 10928 5040 10934 5052
rect 11977 5049 11989 5052
rect 12023 5080 12035 5083
rect 13722 5080 13728 5092
rect 12023 5052 13728 5080
rect 12023 5049 12035 5052
rect 11977 5043 12035 5049
rect 13722 5040 13728 5052
rect 13780 5080 13786 5092
rect 13817 5083 13875 5089
rect 13817 5080 13829 5083
rect 13780 5052 13829 5080
rect 13780 5040 13786 5052
rect 13817 5049 13829 5052
rect 13863 5049 13875 5083
rect 13817 5043 13875 5049
rect 18785 5083 18843 5089
rect 18785 5049 18797 5083
rect 18831 5080 18843 5083
rect 20070 5080 20076 5092
rect 18831 5052 20076 5080
rect 18831 5049 18843 5052
rect 18785 5043 18843 5049
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 20165 5083 20223 5089
rect 20165 5049 20177 5083
rect 20211 5080 20223 5083
rect 22922 5080 22928 5092
rect 20211 5052 22928 5080
rect 20211 5049 20223 5052
rect 20165 5043 20223 5049
rect 22922 5040 22928 5052
rect 22980 5040 22986 5092
rect 23109 5083 23167 5089
rect 23109 5049 23121 5083
rect 23155 5080 23167 5083
rect 23934 5080 23940 5092
rect 23155 5052 23940 5080
rect 23155 5049 23167 5052
rect 23109 5043 23167 5049
rect 23934 5040 23940 5052
rect 23992 5040 23998 5092
rect 24394 5080 24400 5092
rect 24355 5052 24400 5080
rect 24394 5040 24400 5052
rect 24452 5040 24458 5092
rect 6144 4984 7328 5012
rect 7745 5015 7803 5021
rect 6144 4972 6150 4984
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 7834 5012 7840 5024
rect 7791 4984 7840 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 9214 5012 9220 5024
rect 8260 4984 9220 5012
rect 8260 4972 8266 4984
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9456 4984 9781 5012
rect 9456 4972 9462 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 9769 4975 9827 4981
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 9916 4984 10793 5012
rect 9916 4972 9922 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11204 4984 11529 5012
rect 11204 4972 11210 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 16390 5012 16396 5024
rect 11756 4984 16396 5012
rect 11756 4972 11762 4984
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 19426 5012 19432 5024
rect 19387 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20772 4984 20821 5012
rect 20772 4972 20778 4984
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 20809 4975 20867 4981
rect 23569 5015 23627 5021
rect 23569 4981 23581 5015
rect 23615 5012 23627 5015
rect 24412 5012 24440 5040
rect 23615 4984 24440 5012
rect 23615 4981 23627 4984
rect 23569 4975 23627 4981
rect 25406 4972 25412 5024
rect 25464 5012 25470 5024
rect 26786 5012 26792 5024
rect 25464 4984 26792 5012
rect 25464 4972 25470 4984
rect 26786 4972 26792 4984
rect 26844 4972 26850 5024
rect 27080 5012 27108 5188
rect 27246 5176 27252 5188
rect 27304 5176 27310 5228
rect 27516 5219 27574 5225
rect 27516 5185 27528 5219
rect 27562 5216 27574 5219
rect 27562 5188 29224 5216
rect 27562 5185 27574 5188
rect 27516 5179 27574 5185
rect 29196 5148 29224 5188
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 30392 5225 30420 5256
rect 31294 5244 31300 5256
rect 31352 5244 31358 5296
rect 33962 5284 33968 5296
rect 32876 5256 33968 5284
rect 30377 5219 30435 5225
rect 29328 5188 29373 5216
rect 29328 5176 29334 5188
rect 30377 5185 30389 5219
rect 30423 5185 30435 5219
rect 30377 5179 30435 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5216 30619 5219
rect 30650 5216 30656 5228
rect 30607 5188 30656 5216
rect 30607 5185 30619 5188
rect 30561 5179 30619 5185
rect 30650 5176 30656 5188
rect 30708 5176 30714 5228
rect 30834 5216 30840 5228
rect 30795 5188 30840 5216
rect 30834 5176 30840 5188
rect 30892 5176 30898 5228
rect 30926 5176 30932 5228
rect 30984 5216 30990 5228
rect 30984 5188 31029 5216
rect 30984 5176 30990 5188
rect 31110 5176 31116 5228
rect 31168 5216 31174 5228
rect 32876 5225 32904 5256
rect 33962 5244 33968 5256
rect 34020 5244 34026 5296
rect 34057 5287 34115 5293
rect 34057 5253 34069 5287
rect 34103 5284 34115 5287
rect 34790 5284 34796 5296
rect 34103 5256 34796 5284
rect 34103 5253 34115 5256
rect 34057 5247 34115 5253
rect 34790 5244 34796 5256
rect 34848 5244 34854 5296
rect 34968 5287 35026 5293
rect 34968 5253 34980 5287
rect 35014 5284 35026 5287
rect 37182 5284 37188 5296
rect 35014 5256 37188 5284
rect 35014 5253 35026 5256
rect 34968 5247 35026 5253
rect 37182 5244 37188 5256
rect 37240 5244 37246 5296
rect 32769 5219 32827 5225
rect 32769 5216 32781 5219
rect 31168 5188 32781 5216
rect 31168 5176 31174 5188
rect 32769 5185 32781 5188
rect 32815 5185 32827 5219
rect 32769 5179 32827 5185
rect 32861 5219 32919 5225
rect 32861 5185 32873 5219
rect 32907 5185 32919 5219
rect 32861 5179 32919 5185
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5216 33195 5219
rect 33594 5216 33600 5228
rect 33183 5188 33600 5216
rect 33183 5185 33195 5188
rect 33137 5179 33195 5185
rect 33594 5176 33600 5188
rect 33652 5176 33658 5228
rect 33870 5216 33876 5228
rect 33831 5188 33876 5216
rect 33870 5176 33876 5188
rect 33928 5176 33934 5228
rect 34698 5216 34704 5228
rect 34659 5188 34704 5216
rect 34698 5176 34704 5188
rect 34756 5176 34762 5228
rect 35894 5176 35900 5228
rect 35952 5216 35958 5228
rect 36725 5219 36783 5225
rect 36725 5216 36737 5219
rect 35952 5188 36737 5216
rect 35952 5176 35958 5188
rect 36725 5185 36737 5188
rect 36771 5185 36783 5219
rect 37826 5216 37832 5228
rect 37787 5188 37832 5216
rect 36725 5179 36783 5185
rect 37826 5176 37832 5188
rect 37884 5176 37890 5228
rect 31846 5148 31852 5160
rect 29196 5120 31852 5148
rect 31846 5108 31852 5120
rect 31904 5108 31910 5160
rect 32490 5108 32496 5160
rect 32548 5148 32554 5160
rect 33045 5151 33103 5157
rect 33045 5148 33057 5151
rect 32548 5120 33057 5148
rect 32548 5108 32554 5120
rect 33045 5117 33057 5120
rect 33091 5117 33103 5151
rect 33045 5111 33103 5117
rect 28534 5040 28540 5092
rect 28592 5080 28598 5092
rect 30650 5080 30656 5092
rect 28592 5052 30328 5080
rect 30611 5052 30656 5080
rect 28592 5040 28598 5052
rect 27522 5012 27528 5024
rect 27080 4984 27528 5012
rect 27522 4972 27528 4984
rect 27580 4972 27586 5024
rect 29089 5015 29147 5021
rect 29089 4981 29101 5015
rect 29135 5012 29147 5015
rect 30190 5012 30196 5024
rect 29135 4984 30196 5012
rect 29135 4981 29147 4984
rect 29089 4975 29147 4981
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 30300 5012 30328 5052
rect 30650 5040 30656 5052
rect 30708 5040 30714 5092
rect 32585 5083 32643 5089
rect 32585 5049 32597 5083
rect 32631 5080 32643 5083
rect 32858 5080 32864 5092
rect 32631 5052 32864 5080
rect 32631 5049 32643 5052
rect 32585 5043 32643 5049
rect 32858 5040 32864 5052
rect 32916 5080 32922 5092
rect 34514 5080 34520 5092
rect 32916 5052 34520 5080
rect 32916 5040 32922 5052
rect 34514 5040 34520 5052
rect 34572 5040 34578 5092
rect 35434 5012 35440 5024
rect 30300 4984 35440 5012
rect 35434 4972 35440 4984
rect 35492 5012 35498 5024
rect 35802 5012 35808 5024
rect 35492 4984 35808 5012
rect 35492 4972 35498 4984
rect 35802 4972 35808 4984
rect 35860 4972 35866 5024
rect 36541 5015 36599 5021
rect 36541 4981 36553 5015
rect 36587 5012 36599 5015
rect 37826 5012 37832 5024
rect 36587 4984 37832 5012
rect 36587 4981 36599 4984
rect 36541 4975 36599 4981
rect 37826 4972 37832 4984
rect 37884 4972 37890 5024
rect 38013 5015 38071 5021
rect 38013 4981 38025 5015
rect 38059 5012 38071 5015
rect 39758 5012 39764 5024
rect 38059 4984 39764 5012
rect 38059 4981 38071 4984
rect 38013 4975 38071 4981
rect 39758 4972 39764 4984
rect 39816 4972 39822 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5040 4780 8156 4808
rect 5040 4768 5046 4780
rect 4249 4743 4307 4749
rect 4249 4709 4261 4743
rect 4295 4740 4307 4743
rect 5442 4740 5448 4752
rect 4295 4712 5448 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 8128 4740 8156 4780
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8662 4808 8668 4820
rect 8260 4780 8668 4808
rect 8260 4768 8266 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 8996 4780 9781 4808
rect 8996 4768 9002 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10686 4808 10692 4820
rect 10551 4780 10692 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 12066 4808 12072 4820
rect 11020 4780 12072 4808
rect 11020 4768 11026 4780
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12802 4808 12808 4820
rect 12763 4780 12808 4808
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 12952 4780 13584 4808
rect 12952 4768 12958 4780
rect 13556 4752 13584 4780
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 16209 4811 16267 4817
rect 16209 4808 16221 4811
rect 14700 4780 16221 4808
rect 14700 4768 14706 4780
rect 16209 4777 16221 4780
rect 16255 4777 16267 4811
rect 16209 4771 16267 4777
rect 16945 4811 17003 4817
rect 16945 4777 16957 4811
rect 16991 4808 17003 4811
rect 17034 4808 17040 4820
rect 16991 4780 17040 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 20622 4808 20628 4820
rect 18840 4780 20484 4808
rect 20583 4780 20628 4808
rect 18840 4768 18846 4780
rect 10226 4740 10232 4752
rect 8128 4712 10232 4740
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 10410 4700 10416 4752
rect 10468 4740 10474 4752
rect 13538 4740 13544 4752
rect 10468 4712 13400 4740
rect 13499 4712 13544 4740
rect 10468 4700 10474 4712
rect 6822 4672 6828 4684
rect 6012 4644 6684 4672
rect 6783 4644 6828 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3252 4536 3280 4567
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4212 4576 4445 4604
rect 4212 4564 4218 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5166 4604 5172 4616
rect 5123 4576 5172 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6012 4604 6040 4644
rect 5767 4576 6040 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6144 4576 6377 4604
rect 6144 4564 6150 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6656 4604 6684 4644
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 8352 4644 9413 4672
rect 8352 4632 8358 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 10594 4672 10600 4684
rect 9401 4635 9459 4641
rect 9508 4644 10600 4672
rect 6914 4604 6920 4616
rect 6656 4576 6920 4604
rect 6365 4567 6423 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 7098 4613 7104 4616
rect 7092 4604 7104 4613
rect 7059 4576 7104 4604
rect 7092 4567 7104 4576
rect 7098 4564 7104 4567
rect 7156 4564 7162 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 9508 4604 9536 4644
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 13372 4672 13400 4712
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 15930 4700 15936 4752
rect 15988 4740 15994 4752
rect 17865 4743 17923 4749
rect 17865 4740 17877 4743
rect 15988 4712 17877 4740
rect 15988 4700 15994 4712
rect 17865 4709 17877 4712
rect 17911 4709 17923 4743
rect 17865 4703 17923 4709
rect 15562 4672 15568 4684
rect 13044 4644 13308 4672
rect 13372 4644 15568 4672
rect 13044 4632 13050 4644
rect 7432 4576 9536 4604
rect 9585 4607 9643 4613
rect 7432 4564 7438 4576
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 9858 4604 9864 4616
rect 9631 4576 9864 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10376 4576 10425 4604
rect 10376 4564 10382 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 10502 4564 10508 4616
rect 10560 4604 10566 4616
rect 12526 4604 12532 4616
rect 10560 4576 10605 4604
rect 12487 4576 12532 4604
rect 10560 4564 10566 4576
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4604 12679 4607
rect 13170 4604 13176 4616
rect 12667 4576 13176 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 13280 4604 13308 4644
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17313 4675 17371 4681
rect 17313 4672 17325 4675
rect 17092 4644 17325 4672
rect 17092 4632 17098 4644
rect 17313 4641 17325 4644
rect 17359 4641 17371 4675
rect 17313 4635 17371 4641
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4672 17463 4675
rect 18322 4672 18328 4684
rect 17451 4644 18328 4672
rect 17451 4641 17463 4644
rect 17405 4635 17463 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18414 4632 18420 4684
rect 18472 4672 18478 4684
rect 19242 4672 19248 4684
rect 18472 4644 19248 4672
rect 18472 4632 18478 4644
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 20456 4672 20484 4780
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 23842 4808 23848 4820
rect 23803 4780 23848 4808
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 26418 4808 26424 4820
rect 24688 4780 26424 4808
rect 22462 4672 22468 4684
rect 20456 4644 22094 4672
rect 22423 4644 22468 4672
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13280 4576 14473 4604
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4604 14979 4607
rect 15010 4604 15016 4616
rect 14967 4576 15016 4604
rect 14967 4573 14979 4576
rect 14921 4567 14979 4573
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 15286 4604 15292 4616
rect 15243 4576 15292 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 16390 4604 16396 4616
rect 16351 4576 16396 4604
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 19058 4604 19064 4616
rect 18739 4576 19064 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 5350 4536 5356 4548
rect 3252 4508 5356 4536
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 10226 4536 10232 4548
rect 5552 4508 10088 4536
rect 10187 4508 10232 4536
rect 1397 4471 1455 4477
rect 1397 4437 1409 4471
rect 1443 4468 1455 4471
rect 1854 4468 1860 4480
rect 1443 4440 1860 4468
rect 1443 4437 1455 4440
rect 1397 4431 1455 4437
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4890 4468 4896 4480
rect 4851 4440 4896 4468
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5552 4477 5580 4508
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4437 5595 4471
rect 5537 4431 5595 4437
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 8754 4468 8760 4480
rect 6227 4440 8760 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 10060 4468 10088 4508
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 10962 4536 10968 4548
rect 10612 4508 10968 4536
rect 10612 4468 10640 4508
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11146 4536 11152 4548
rect 11107 4508 11152 4536
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11333 4539 11391 4545
rect 11333 4505 11345 4539
rect 11379 4536 11391 4539
rect 11606 4536 11612 4548
rect 11379 4508 11612 4536
rect 11379 4505 11391 4508
rect 11333 4499 11391 4505
rect 10060 4440 10640 4468
rect 10689 4471 10747 4477
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 10778 4468 10784 4480
rect 10735 4440 10784 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11348 4468 11376 4499
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 11790 4496 11796 4548
rect 11848 4536 11854 4548
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 11848 4508 12357 4536
rect 11848 4496 11854 4508
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 12345 4499 12403 4505
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 13357 4539 13415 4545
rect 13357 4536 13369 4539
rect 12768 4508 13369 4536
rect 12768 4496 12774 4508
rect 13357 4505 13369 4508
rect 13403 4505 13415 4539
rect 13357 4499 13415 4505
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 18064 4536 18092 4567
rect 16540 4508 18092 4536
rect 18524 4536 18552 4567
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19512 4607 19570 4613
rect 19512 4573 19524 4607
rect 19558 4604 19570 4607
rect 19978 4604 19984 4616
rect 19558 4576 19984 4604
rect 19558 4573 19570 4576
rect 19512 4567 19570 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 21082 4604 21088 4616
rect 20864 4576 21088 4604
rect 20864 4564 20870 4576
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 22066 4604 22094 4644
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 22554 4604 22560 4616
rect 22066 4576 22560 4604
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23072 4576 23520 4604
rect 23072 4564 23078 4576
rect 20438 4536 20444 4548
rect 18524 4508 20444 4536
rect 16540 4496 16546 4508
rect 20438 4496 20444 4508
rect 20496 4496 20502 4548
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 21269 4539 21327 4545
rect 21269 4536 21281 4539
rect 21048 4508 21281 4536
rect 21048 4496 21054 4508
rect 21269 4505 21281 4508
rect 21315 4505 21327 4539
rect 22732 4539 22790 4545
rect 21269 4499 21327 4505
rect 21376 4508 22094 4536
rect 11112 4440 11376 4468
rect 11517 4471 11575 4477
rect 11112 4428 11118 4440
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 13446 4468 13452 4480
rect 11563 4440 13452 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14274 4468 14280 4480
rect 14235 4440 14280 4468
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 19978 4468 19984 4480
rect 18647 4440 19984 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 21376 4468 21404 4508
rect 20220 4440 21404 4468
rect 21453 4471 21511 4477
rect 20220 4428 20226 4440
rect 21453 4437 21465 4471
rect 21499 4468 21511 4471
rect 21818 4468 21824 4480
rect 21499 4440 21824 4468
rect 21499 4437 21511 4440
rect 21453 4431 21511 4437
rect 21818 4428 21824 4440
rect 21876 4428 21882 4480
rect 22066 4468 22094 4508
rect 22732 4505 22744 4539
rect 22778 4536 22790 4539
rect 23382 4536 23388 4548
rect 22778 4508 23388 4536
rect 22778 4505 22790 4508
rect 22732 4499 22790 4505
rect 23382 4496 23388 4508
rect 23440 4496 23446 4548
rect 23492 4536 23520 4576
rect 23934 4564 23940 4616
rect 23992 4604 23998 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23992 4576 24593 4604
rect 23992 4564 23998 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 24397 4539 24455 4545
rect 24397 4536 24409 4539
rect 23492 4508 24409 4536
rect 24397 4505 24409 4508
rect 24443 4505 24455 4539
rect 24397 4499 24455 4505
rect 24688 4468 24716 4780
rect 26418 4768 26424 4780
rect 26476 4768 26482 4820
rect 26694 4808 26700 4820
rect 26655 4780 26700 4808
rect 26694 4768 26700 4780
rect 26752 4768 26758 4820
rect 26786 4768 26792 4820
rect 26844 4808 26850 4820
rect 28074 4808 28080 4820
rect 26844 4780 28080 4808
rect 26844 4768 26850 4780
rect 28074 4768 28080 4780
rect 28132 4768 28138 4820
rect 28169 4811 28227 4817
rect 28169 4777 28181 4811
rect 28215 4808 28227 4811
rect 29454 4808 29460 4820
rect 28215 4780 29460 4808
rect 28215 4777 28227 4780
rect 28169 4771 28227 4777
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 29638 4768 29644 4820
rect 29696 4808 29702 4820
rect 31110 4808 31116 4820
rect 29696 4780 31116 4808
rect 29696 4768 29702 4780
rect 31110 4768 31116 4780
rect 31168 4768 31174 4820
rect 33134 4808 33140 4820
rect 31726 4780 33140 4808
rect 26237 4743 26295 4749
rect 26237 4709 26249 4743
rect 26283 4740 26295 4743
rect 31726 4740 31754 4780
rect 33134 4768 33140 4780
rect 33192 4768 33198 4820
rect 33594 4808 33600 4820
rect 33555 4780 33600 4808
rect 33594 4768 33600 4780
rect 33652 4768 33658 4820
rect 35161 4811 35219 4817
rect 35161 4777 35173 4811
rect 35207 4808 35219 4811
rect 37366 4808 37372 4820
rect 35207 4780 37372 4808
rect 35207 4777 35219 4780
rect 35161 4771 35219 4777
rect 37366 4768 37372 4780
rect 37424 4768 37430 4820
rect 26283 4712 31754 4740
rect 36265 4743 36323 4749
rect 26283 4709 26295 4712
rect 26237 4703 26295 4709
rect 36265 4709 36277 4743
rect 36311 4740 36323 4743
rect 37274 4740 37280 4752
rect 36311 4712 37280 4740
rect 36311 4709 36323 4712
rect 36265 4703 36323 4709
rect 37274 4700 37280 4712
rect 37332 4700 37338 4752
rect 24765 4675 24823 4681
rect 24765 4641 24777 4675
rect 24811 4672 24823 4675
rect 27706 4672 27712 4684
rect 24811 4644 27712 4672
rect 24811 4641 24823 4644
rect 24765 4635 24823 4641
rect 27706 4632 27712 4644
rect 27764 4632 27770 4684
rect 28074 4632 28080 4684
rect 28132 4672 28138 4684
rect 28132 4644 29776 4672
rect 28132 4632 28138 4644
rect 25406 4604 25412 4616
rect 25367 4576 25412 4604
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 26881 4607 26939 4613
rect 26881 4604 26893 4607
rect 25516 4576 26893 4604
rect 24854 4496 24860 4548
rect 24912 4536 24918 4548
rect 25516 4536 25544 4576
rect 26881 4573 26893 4576
rect 26927 4573 26939 4607
rect 26881 4567 26939 4573
rect 27522 4564 27528 4616
rect 27580 4604 27586 4616
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27580 4576 27813 4604
rect 27580 4564 27586 4576
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 27985 4607 28043 4613
rect 27985 4573 27997 4607
rect 28031 4604 28043 4607
rect 28350 4604 28356 4616
rect 28031 4576 28356 4604
rect 28031 4573 28043 4576
rect 27985 4567 28043 4573
rect 28350 4564 28356 4576
rect 28408 4564 28414 4616
rect 28626 4604 28632 4616
rect 28587 4576 28632 4604
rect 28626 4564 28632 4576
rect 28684 4564 28690 4616
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 28994 4604 29000 4616
rect 28859 4576 29000 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 29748 4613 29776 4644
rect 29822 4632 29828 4684
rect 29880 4672 29886 4684
rect 36906 4672 36912 4684
rect 29880 4644 31064 4672
rect 29880 4632 29886 4644
rect 31036 4613 31064 4644
rect 34900 4644 36912 4672
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 30377 4607 30435 4613
rect 30377 4573 30389 4607
rect 30423 4573 30435 4607
rect 30377 4567 30435 4573
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4573 31079 4607
rect 31478 4604 31484 4616
rect 31439 4576 31484 4604
rect 31021 4567 31079 4573
rect 24912 4508 25544 4536
rect 25869 4539 25927 4545
rect 24912 4496 24918 4508
rect 25869 4505 25881 4539
rect 25915 4505 25927 4539
rect 26050 4536 26056 4548
rect 26011 4508 26056 4536
rect 25869 4499 25927 4505
rect 22066 4440 24716 4468
rect 25130 4428 25136 4480
rect 25188 4468 25194 4480
rect 25225 4471 25283 4477
rect 25225 4468 25237 4471
rect 25188 4440 25237 4468
rect 25188 4428 25194 4440
rect 25225 4437 25237 4440
rect 25271 4437 25283 4471
rect 25884 4468 25912 4499
rect 26050 4496 26056 4508
rect 26108 4496 26114 4548
rect 28258 4496 28264 4548
rect 28316 4536 28322 4548
rect 30392 4536 30420 4567
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 31665 4607 31723 4613
rect 31665 4573 31677 4607
rect 31711 4573 31723 4607
rect 32214 4604 32220 4616
rect 32175 4576 32220 4604
rect 31665 4567 31723 4573
rect 31680 4536 31708 4567
rect 32214 4564 32220 4576
rect 32272 4564 32278 4616
rect 32484 4607 32542 4613
rect 32484 4573 32496 4607
rect 32530 4604 32542 4607
rect 34900 4604 34928 4644
rect 36906 4632 36912 4644
rect 36964 4632 36970 4684
rect 32530 4576 34928 4604
rect 34977 4607 35035 4613
rect 32530 4573 32542 4576
rect 32484 4567 32542 4573
rect 34977 4573 34989 4607
rect 35023 4604 35035 4607
rect 35710 4604 35716 4616
rect 35023 4576 35716 4604
rect 35023 4573 35035 4576
rect 34977 4567 35035 4573
rect 35710 4564 35716 4576
rect 35768 4564 35774 4616
rect 35802 4564 35808 4616
rect 35860 4604 35866 4616
rect 36446 4604 36452 4616
rect 35860 4576 35905 4604
rect 36407 4576 36452 4604
rect 35860 4564 35866 4576
rect 36446 4564 36452 4576
rect 36504 4564 36510 4616
rect 36538 4564 36544 4616
rect 36596 4604 36602 4616
rect 37369 4607 37427 4613
rect 37369 4604 37381 4607
rect 36596 4576 37381 4604
rect 36596 4564 36602 4576
rect 37369 4573 37381 4576
rect 37415 4573 37427 4607
rect 37826 4604 37832 4616
rect 37787 4576 37832 4604
rect 37369 4567 37427 4573
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 28316 4508 30420 4536
rect 30760 4508 31754 4536
rect 28316 4496 28322 4508
rect 27522 4468 27528 4480
rect 25884 4440 27528 4468
rect 25225 4431 25283 4437
rect 27522 4428 27528 4440
rect 27580 4428 27586 4480
rect 28442 4428 28448 4480
rect 28500 4468 28506 4480
rect 28721 4471 28779 4477
rect 28721 4468 28733 4471
rect 28500 4440 28733 4468
rect 28500 4428 28506 4440
rect 28721 4437 28733 4440
rect 28767 4437 28779 4471
rect 29546 4468 29552 4480
rect 29507 4440 29552 4468
rect 28721 4431 28779 4437
rect 29546 4428 29552 4440
rect 29604 4428 29610 4480
rect 29730 4428 29736 4480
rect 29788 4468 29794 4480
rect 30193 4471 30251 4477
rect 30193 4468 30205 4471
rect 29788 4440 30205 4468
rect 29788 4428 29794 4440
rect 30193 4437 30205 4440
rect 30239 4437 30251 4471
rect 30193 4431 30251 4437
rect 30282 4428 30288 4480
rect 30340 4468 30346 4480
rect 30760 4468 30788 4508
rect 30340 4440 30788 4468
rect 30837 4471 30895 4477
rect 30340 4428 30346 4440
rect 30837 4437 30849 4471
rect 30883 4468 30895 4471
rect 31018 4468 31024 4480
rect 30883 4440 31024 4468
rect 30883 4437 30895 4440
rect 30837 4431 30895 4437
rect 31018 4428 31024 4440
rect 31076 4428 31082 4480
rect 31570 4468 31576 4480
rect 31531 4440 31576 4468
rect 31570 4428 31576 4440
rect 31628 4428 31634 4480
rect 31726 4468 31754 4508
rect 33870 4496 33876 4548
rect 33928 4536 33934 4548
rect 34793 4539 34851 4545
rect 34793 4536 34805 4539
rect 33928 4508 34805 4536
rect 33928 4496 33934 4508
rect 34793 4505 34805 4508
rect 34839 4536 34851 4539
rect 36262 4536 36268 4548
rect 34839 4508 36268 4536
rect 34839 4505 34851 4508
rect 34793 4499 34851 4505
rect 36262 4496 36268 4508
rect 36320 4496 36326 4548
rect 32306 4468 32312 4480
rect 31726 4440 32312 4468
rect 32306 4428 32312 4440
rect 32364 4428 32370 4480
rect 35618 4468 35624 4480
rect 35579 4440 35624 4468
rect 35618 4428 35624 4440
rect 35676 4428 35682 4480
rect 37185 4471 37243 4477
rect 37185 4437 37197 4471
rect 37231 4468 37243 4471
rect 37826 4468 37832 4480
rect 37231 4440 37832 4468
rect 37231 4437 37243 4440
rect 37185 4431 37243 4437
rect 37826 4428 37832 4440
rect 37884 4428 37890 4480
rect 38013 4471 38071 4477
rect 38013 4437 38025 4471
rect 38059 4468 38071 4471
rect 39022 4468 39028 4480
rect 38059 4440 39028 4468
rect 38059 4437 38071 4440
rect 38013 4431 38071 4437
rect 39022 4428 39028 4440
rect 39080 4428 39086 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3421 4267 3479 4273
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 5626 4264 5632 4276
rect 3467 4236 5304 4264
rect 5587 4236 5632 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 992 4100 1593 4128
rect 992 4088 998 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 3053 4131 3111 4137
rect 2639 4100 2774 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2746 4060 2774 4100
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3602 4128 3608 4140
rect 3099 4100 3608 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3896 4137 3924 4236
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5276 4196 5304 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 5736 4236 7954 4264
rect 5736 4196 5764 4236
rect 7098 4196 7104 4208
rect 5132 4168 5212 4196
rect 5276 4168 5764 4196
rect 7059 4168 7104 4196
rect 5132 4156 5138 4168
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 5184 4137 5212 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 5169 4131 5227 4137
rect 4580 4100 4625 4128
rect 4580 4088 4586 4100
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6730 4128 6736 4140
rect 5859 4100 6736 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7708 4100 7757 4128
rect 7708 4088 7714 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 4706 4060 4712 4072
rect 2746 4032 4712 4060
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 7834 4060 7840 4072
rect 7795 4032 7840 4060
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 7926 4060 7954 4236
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 9628 4264 9634 4276
rect 8904 4236 9634 4264
rect 8904 4224 8910 4236
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8202 4128 8208 4140
rect 8067 4100 8208 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9306 4128 9312 4140
rect 8987 4100 9312 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9508 4128 9536 4236
rect 9628 4224 9634 4236
rect 9686 4224 9692 4276
rect 13722 4264 13728 4276
rect 12820 4236 13728 4264
rect 11977 4199 12035 4205
rect 11977 4165 11989 4199
rect 12023 4196 12035 4199
rect 12710 4196 12716 4208
rect 12023 4168 12716 4196
rect 12023 4165 12035 4168
rect 11977 4159 12035 4165
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 12820 4205 12848 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 20162 4264 20168 4276
rect 16448 4236 20168 4264
rect 16448 4224 16454 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 21177 4267 21235 4273
rect 21177 4233 21189 4267
rect 21223 4264 21235 4267
rect 22646 4264 22652 4276
rect 21223 4236 22652 4264
rect 21223 4233 21235 4236
rect 21177 4227 21235 4233
rect 22646 4224 22652 4236
rect 22704 4264 22710 4276
rect 25406 4264 25412 4276
rect 22704 4236 25412 4264
rect 22704 4224 22710 4236
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 25869 4267 25927 4273
rect 25869 4233 25881 4267
rect 25915 4264 25927 4267
rect 26050 4264 26056 4276
rect 25915 4236 26056 4264
rect 25915 4233 25927 4236
rect 25869 4227 25927 4233
rect 12805 4199 12863 4205
rect 12805 4165 12817 4199
rect 12851 4165 12863 4199
rect 15286 4196 15292 4208
rect 12805 4159 12863 4165
rect 13740 4168 15292 4196
rect 9568 4131 9626 4137
rect 9568 4128 9580 4131
rect 9508 4100 9580 4128
rect 9568 4097 9580 4100
rect 9614 4097 9626 4131
rect 9568 4091 9626 4097
rect 9674 4088 9680 4140
rect 9732 4137 9738 4140
rect 9732 4131 9765 4137
rect 9753 4097 9765 4131
rect 9732 4091 9765 4097
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 9732 4088 9738 4091
rect 9214 4060 9220 4072
rect 7926 4032 9220 4060
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9968 4060 9996 4091
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10100 4100 10609 4128
rect 10100 4088 10106 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10965 4131 11023 4137
rect 10744 4100 10789 4128
rect 10744 4088 10750 4100
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 12158 4128 12164 4140
rect 12119 4100 12164 4128
rect 10965 4091 11023 4097
rect 10870 4060 10876 4072
rect 9600 4032 9996 4060
rect 10831 4032 10876 4060
rect 2406 3992 2412 4004
rect 2367 3964 2412 3992
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 2866 3992 2872 4004
rect 2827 3964 2872 3992
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 9600 3992 9628 4032
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 3108 3964 9628 3992
rect 9861 3995 9919 4001
rect 3108 3952 3114 3964
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 10042 3992 10048 4004
rect 9907 3964 10048 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 10980 3992 11008 4091
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12618 4128 12624 4140
rect 12579 4100 12624 4128
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12905 4131 12963 4137
rect 12905 4097 12917 4131
rect 12951 4097 12963 4131
rect 12905 4091 12963 4097
rect 13035 4131 13093 4137
rect 13035 4097 13047 4131
rect 13081 4128 13093 4131
rect 13740 4128 13768 4168
rect 15286 4156 15292 4168
rect 15344 4196 15350 4208
rect 19058 4196 19064 4208
rect 15344 4168 17080 4196
rect 15344 4156 15350 4168
rect 13081 4100 13768 4128
rect 13817 4131 13875 4137
rect 13081 4097 13093 4100
rect 13035 4091 13093 4097
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 14182 4128 14188 4140
rect 13863 4100 14188 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 12913 4060 12941 4091
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 16114 4128 16120 4140
rect 16075 4100 16120 4128
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16758 4128 16764 4140
rect 16715 4100 16764 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17052 4137 17080 4168
rect 18524 4168 19064 4196
rect 18524 4137 18552 4168
rect 19058 4156 19064 4168
rect 19116 4196 19122 4208
rect 20990 4196 20996 4208
rect 19116 4168 19380 4196
rect 19116 4156 19122 4168
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 16941 4131 16999 4137
rect 16941 4097 16953 4131
rect 16987 4097 16999 4131
rect 16941 4091 16999 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 18874 4128 18880 4140
rect 18739 4100 18880 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 11480 4032 12941 4060
rect 13633 4063 13691 4069
rect 11480 4020 11486 4032
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14274 4060 14280 4072
rect 13679 4032 14280 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 15102 4060 15108 4072
rect 14967 4032 15108 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 10652 3964 11008 3992
rect 10652 3952 10658 3964
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 14660 3992 14688 4023
rect 15102 4020 15108 4032
rect 15160 4060 15166 4072
rect 16868 4060 16896 4091
rect 15160 4032 16896 4060
rect 15160 4020 15166 4032
rect 15010 3992 15016 4004
rect 11204 3964 14136 3992
rect 14660 3964 15016 3992
rect 11204 3952 11210 3964
rect 1397 3927 1455 3933
rect 1397 3893 1409 3927
rect 1443 3924 1455 3927
rect 2038 3924 2044 3936
rect 1443 3896 2044 3924
rect 1443 3893 1455 3896
rect 1397 3887 1455 3893
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4614 3924 4620 3936
rect 4387 3896 4620 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 7285 3927 7343 3933
rect 7285 3924 7297 3927
rect 5868 3896 7297 3924
rect 5868 3884 5874 3896
rect 7285 3893 7297 3896
rect 7331 3893 7343 3927
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7285 3887 7343 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7984 3896 8217 3924
rect 7984 3884 7990 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9030 3924 9036 3936
rect 8803 3896 9036 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9398 3924 9404 3936
rect 9359 3896 9404 3924
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12952 3896 13185 3924
rect 12952 3884 12958 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13998 3924 14004 3936
rect 13959 3896 14004 3924
rect 13173 3887 13231 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14108 3924 14136 3964
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 16951 3992 16979 4091
rect 18064 4060 18092 4091
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19352 4137 19380 4168
rect 20916 4168 20996 4196
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4097 19395 4131
rect 19337 4091 19395 4097
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20916 4137 20944 4168
rect 20990 4156 20996 4168
rect 21048 4156 21054 4208
rect 22741 4199 22799 4205
rect 22741 4196 22753 4199
rect 22112 4168 22753 4196
rect 22112 4140 22140 4168
rect 22741 4165 22753 4168
rect 22787 4165 22799 4199
rect 25774 4196 25780 4208
rect 22741 4159 22799 4165
rect 22940 4168 25780 4196
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 20128 4100 20177 4128
rect 20128 4088 20134 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 20901 4131 20959 4137
rect 20901 4097 20913 4131
rect 20947 4097 20959 4131
rect 21082 4128 21088 4140
rect 21043 4100 21088 4128
rect 20901 4091 20959 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 21634 4088 21640 4140
rect 21692 4128 21698 4140
rect 22005 4131 22063 4137
rect 21692 4100 21956 4128
rect 21692 4088 21698 4100
rect 21542 4060 21548 4072
rect 18064 4032 21548 4060
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 21821 4063 21879 4069
rect 21821 4029 21833 4063
rect 21867 4029 21879 4063
rect 21928 4060 21956 4100
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22940 4137 22968 4168
rect 25774 4156 25780 4168
rect 25832 4156 25838 4208
rect 22925 4131 22983 4137
rect 22244 4100 22289 4128
rect 22244 4088 22250 4100
rect 22925 4097 22937 4131
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 23293 4131 23351 4137
rect 23293 4097 23305 4131
rect 23339 4128 23351 4131
rect 23474 4128 23480 4140
rect 23339 4100 23480 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 23032 4060 23060 4091
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 23934 4128 23940 4140
rect 23895 4100 23940 4128
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 24121 4131 24179 4137
rect 24121 4097 24133 4131
rect 24167 4128 24179 4131
rect 24854 4128 24860 4140
rect 24167 4100 24860 4128
rect 24167 4097 24179 4100
rect 24121 4091 24179 4097
rect 24854 4088 24860 4100
rect 24912 4088 24918 4140
rect 25225 4131 25283 4137
rect 25225 4097 25237 4131
rect 25271 4128 25283 4131
rect 25884 4128 25912 4227
rect 26050 4224 26056 4236
rect 26108 4224 26114 4276
rect 27522 4264 27528 4276
rect 26988 4236 27528 4264
rect 26988 4205 27016 4236
rect 27522 4224 27528 4236
rect 27580 4224 27586 4276
rect 28718 4264 28724 4276
rect 27724 4236 28724 4264
rect 26973 4199 27031 4205
rect 26973 4165 26985 4199
rect 27019 4165 27031 4199
rect 26973 4159 27031 4165
rect 27157 4199 27215 4205
rect 27157 4165 27169 4199
rect 27203 4196 27215 4199
rect 27724 4196 27752 4236
rect 28718 4224 28724 4236
rect 28776 4224 28782 4276
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 29052 4236 29960 4264
rect 29052 4224 29058 4236
rect 28810 4196 28816 4208
rect 27203 4168 27752 4196
rect 27816 4168 28816 4196
rect 27203 4165 27215 4168
rect 27157 4159 27215 4165
rect 27816 4140 27844 4168
rect 28810 4156 28816 4168
rect 28868 4156 28874 4208
rect 29638 4196 29644 4208
rect 28903 4168 29644 4196
rect 28903 4140 28931 4168
rect 29638 4156 29644 4168
rect 29696 4156 29702 4208
rect 25271 4100 25912 4128
rect 25271 4097 25283 4100
rect 25225 4091 25283 4097
rect 25958 4088 25964 4140
rect 26016 4128 26022 4140
rect 26053 4131 26111 4137
rect 26053 4128 26065 4131
rect 26016 4100 26065 4128
rect 26016 4088 26022 4100
rect 26053 4097 26065 4100
rect 26099 4097 26111 4131
rect 26053 4091 26111 4097
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 26421 4131 26479 4137
rect 26200 4100 26245 4128
rect 26200 4088 26206 4100
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 26786 4128 26792 4140
rect 26467 4100 26792 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 26786 4088 26792 4100
rect 26844 4088 26850 4140
rect 27338 4128 27344 4140
rect 27299 4100 27344 4128
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 27798 4128 27804 4140
rect 27759 4100 27804 4128
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 27982 4128 27988 4140
rect 27943 4100 27988 4128
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 28169 4131 28227 4137
rect 28169 4097 28181 4131
rect 28215 4128 28227 4131
rect 28258 4128 28264 4140
rect 28215 4100 28264 4128
rect 28215 4097 28227 4100
rect 28169 4091 28227 4097
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 28902 4128 28908 4140
rect 28863 4100 28908 4128
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 28997 4131 29055 4137
rect 28997 4097 29009 4131
rect 29043 4128 29055 4131
rect 29086 4128 29092 4140
rect 29043 4100 29092 4128
rect 29043 4097 29055 4100
rect 28997 4091 29055 4097
rect 29086 4088 29092 4100
rect 29144 4088 29150 4140
rect 29270 4128 29276 4140
rect 29231 4100 29276 4128
rect 29270 4088 29276 4100
rect 29328 4088 29334 4140
rect 29932 4137 29960 4236
rect 35618 4196 35624 4208
rect 30852 4168 32352 4196
rect 30852 4140 30880 4168
rect 32324 4140 32352 4168
rect 34992 4168 35624 4196
rect 29917 4131 29975 4137
rect 29917 4097 29929 4131
rect 29963 4097 29975 4131
rect 29917 4091 29975 4097
rect 30653 4131 30711 4137
rect 30653 4097 30665 4131
rect 30699 4130 30711 4131
rect 30742 4130 30748 4140
rect 30699 4102 30748 4130
rect 30699 4097 30711 4102
rect 30653 4091 30711 4097
rect 30742 4088 30748 4102
rect 30800 4088 30806 4140
rect 30834 4088 30840 4140
rect 30892 4128 30898 4140
rect 31205 4131 31263 4137
rect 30892 4100 30985 4128
rect 30892 4088 30898 4100
rect 31205 4097 31217 4131
rect 31251 4128 31263 4131
rect 31294 4128 31300 4140
rect 31251 4100 31300 4128
rect 31251 4097 31263 4100
rect 31205 4091 31263 4097
rect 31294 4088 31300 4100
rect 31352 4088 31358 4140
rect 32122 4128 32128 4140
rect 32083 4100 32128 4128
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 32306 4128 32312 4140
rect 32219 4100 32312 4128
rect 32306 4088 32312 4100
rect 32364 4088 32370 4140
rect 32401 4131 32459 4137
rect 32401 4097 32413 4131
rect 32447 4128 32459 4131
rect 32582 4128 32588 4140
rect 32447 4100 32588 4128
rect 32447 4097 32459 4100
rect 32401 4091 32459 4097
rect 32582 4088 32588 4100
rect 32640 4088 32646 4140
rect 32677 4131 32735 4137
rect 32677 4097 32689 4131
rect 32723 4128 32735 4131
rect 33134 4128 33140 4140
rect 32723 4100 33140 4128
rect 32723 4097 32735 4100
rect 32677 4091 32735 4097
rect 33134 4088 33140 4100
rect 33192 4088 33198 4140
rect 33502 4128 33508 4140
rect 33463 4100 33508 4128
rect 33502 4088 33508 4100
rect 33560 4088 33566 4140
rect 33965 4131 34023 4137
rect 33965 4097 33977 4131
rect 34011 4128 34023 4131
rect 34054 4128 34060 4140
rect 34011 4100 34060 4128
rect 34011 4097 34023 4100
rect 33965 4091 34023 4097
rect 34054 4088 34060 4100
rect 34112 4088 34118 4140
rect 34992 4137 35020 4168
rect 35618 4156 35624 4168
rect 35676 4156 35682 4208
rect 34149 4131 34207 4137
rect 34149 4097 34161 4131
rect 34195 4097 34207 4131
rect 34149 4091 34207 4097
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4097 35035 4131
rect 34977 4091 35035 4097
rect 21928 4032 23060 4060
rect 21821 4023 21879 4029
rect 15120 3964 16979 3992
rect 15120 3924 15148 3964
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 18012 3964 18521 3992
rect 18012 3952 18018 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 21836 3992 21864 4023
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 23256 4032 23765 4060
rect 23256 4020 23262 4032
rect 23753 4029 23765 4032
rect 23799 4060 23811 4063
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 23799 4032 25053 4060
rect 23799 4029 23811 4032
rect 23753 4023 23811 4029
rect 25041 4029 25053 4032
rect 25087 4060 25099 4063
rect 25130 4060 25136 4072
rect 25087 4032 25136 4060
rect 25087 4029 25099 4032
rect 25041 4023 25099 4029
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25774 4020 25780 4072
rect 25832 4060 25838 4072
rect 30852 4060 30880 4088
rect 25832 4032 29316 4060
rect 25832 4020 25838 4032
rect 22186 3992 22192 4004
rect 21836 3964 22192 3992
rect 18509 3955 18567 3961
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 25409 3995 25467 4001
rect 25409 3961 25421 3995
rect 25455 3992 25467 3995
rect 28994 3992 29000 4004
rect 25455 3964 29000 3992
rect 25455 3961 25467 3964
rect 25409 3955 25467 3961
rect 28994 3952 29000 3964
rect 29052 3952 29058 4004
rect 14108 3896 15148 3924
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 16482 3924 16488 3936
rect 15979 3896 16488 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 16908 3896 17233 3924
rect 16908 3884 16914 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 17865 3927 17923 3933
rect 17865 3893 17877 3927
rect 17911 3924 17923 3927
rect 18230 3924 18236 3936
rect 17911 3896 18236 3924
rect 17911 3893 17923 3896
rect 17865 3887 17923 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 19150 3924 19156 3936
rect 19111 3896 19156 3924
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 20349 3927 20407 3933
rect 20349 3893 20361 3927
rect 20395 3924 20407 3927
rect 22554 3924 22560 3936
rect 20395 3896 22560 3924
rect 20395 3893 20407 3896
rect 20349 3887 20407 3893
rect 22554 3884 22560 3896
rect 22612 3884 22618 3936
rect 23201 3927 23259 3933
rect 23201 3893 23213 3927
rect 23247 3924 23259 3927
rect 24394 3924 24400 3936
rect 23247 3896 24400 3924
rect 23247 3893 23259 3896
rect 23201 3887 23259 3893
rect 24394 3884 24400 3896
rect 24452 3924 24458 3936
rect 26329 3927 26387 3933
rect 26329 3924 26341 3927
rect 24452 3896 26341 3924
rect 24452 3884 24458 3896
rect 26329 3893 26341 3896
rect 26375 3924 26387 3927
rect 28626 3924 28632 3936
rect 26375 3896 28632 3924
rect 26375 3893 26387 3896
rect 26329 3887 26387 3893
rect 28626 3884 28632 3896
rect 28684 3924 28690 3936
rect 29181 3927 29239 3933
rect 29181 3924 29193 3927
rect 28684 3896 29193 3924
rect 28684 3884 28690 3896
rect 29181 3893 29193 3896
rect 29227 3893 29239 3927
rect 29288 3924 29316 4032
rect 29564 4032 30880 4060
rect 30929 4063 30987 4069
rect 29564 3924 29592 4032
rect 30929 4029 30941 4063
rect 30975 4029 30987 4063
rect 30929 4023 30987 4029
rect 31021 4063 31079 4069
rect 31021 4029 31033 4063
rect 31067 4060 31079 4063
rect 32493 4063 32551 4069
rect 31067 4032 31248 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 30834 3952 30840 4004
rect 30892 3992 30898 4004
rect 30944 3992 30972 4023
rect 31220 4004 31248 4032
rect 32493 4029 32505 4063
rect 32539 4060 32551 4063
rect 32950 4060 32956 4072
rect 32539 4032 32956 4060
rect 32539 4029 32551 4032
rect 32493 4023 32551 4029
rect 31110 3992 31116 4004
rect 30892 3964 31116 3992
rect 30892 3952 30898 3964
rect 31110 3952 31116 3964
rect 31168 3952 31174 4004
rect 31202 3952 31208 4004
rect 31260 3992 31266 4004
rect 32508 3992 32536 4023
rect 32950 4020 32956 4032
rect 33008 4020 33014 4072
rect 34164 3992 34192 4091
rect 35066 4088 35072 4140
rect 35124 4128 35130 4140
rect 35713 4131 35771 4137
rect 35124 4100 35169 4128
rect 35124 4088 35130 4100
rect 35713 4097 35725 4131
rect 35759 4128 35771 4131
rect 36630 4128 36636 4140
rect 35759 4100 36492 4128
rect 36591 4100 36636 4128
rect 35759 4097 35771 4100
rect 35713 4091 35771 4097
rect 35253 4063 35311 4069
rect 35253 4029 35265 4063
rect 35299 4060 35311 4063
rect 35894 4060 35900 4072
rect 35299 4032 35900 4060
rect 35299 4029 35311 4032
rect 35253 4023 35311 4029
rect 35894 4020 35900 4032
rect 35952 4020 35958 4072
rect 36464 4001 36492 4100
rect 36630 4088 36636 4100
rect 36688 4088 36694 4140
rect 37826 4128 37832 4140
rect 37787 4100 37832 4128
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 31260 3964 32536 3992
rect 32600 3964 34192 3992
rect 36449 3995 36507 4001
rect 31260 3952 31266 3964
rect 29288 3896 29592 3924
rect 29181 3887 29239 3893
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 29733 3927 29791 3933
rect 29733 3924 29745 3927
rect 29696 3896 29745 3924
rect 29696 3884 29702 3896
rect 29733 3893 29745 3896
rect 29779 3893 29791 3927
rect 31386 3924 31392 3936
rect 31347 3896 31392 3924
rect 29733 3887 29791 3893
rect 31386 3884 31392 3896
rect 31444 3884 31450 3936
rect 32490 3884 32496 3936
rect 32548 3924 32554 3936
rect 32600 3924 32628 3964
rect 36449 3961 36461 3995
rect 36495 3961 36507 3995
rect 36449 3955 36507 3961
rect 32548 3896 32628 3924
rect 32548 3884 32554 3896
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 32861 3927 32919 3933
rect 32861 3924 32873 3927
rect 32732 3896 32873 3924
rect 32732 3884 32738 3896
rect 32861 3893 32873 3896
rect 32907 3893 32919 3927
rect 32861 3887 32919 3893
rect 33321 3927 33379 3933
rect 33321 3893 33333 3927
rect 33367 3924 33379 3927
rect 33870 3924 33876 3936
rect 33367 3896 33876 3924
rect 33367 3893 33379 3896
rect 33321 3887 33379 3893
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 33965 3927 34023 3933
rect 33965 3893 33977 3927
rect 34011 3924 34023 3927
rect 34606 3924 34612 3936
rect 34011 3896 34612 3924
rect 34011 3893 34023 3896
rect 33965 3887 34023 3893
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35897 3927 35955 3933
rect 35897 3924 35909 3927
rect 35400 3896 35909 3924
rect 35400 3884 35406 3896
rect 35897 3893 35909 3896
rect 35943 3893 35955 3927
rect 35897 3887 35955 3893
rect 38013 3927 38071 3933
rect 38013 3893 38025 3927
rect 38059 3924 38071 3927
rect 38286 3924 38292 3936
rect 38059 3896 38292 3924
rect 38059 3893 38071 3896
rect 38013 3887 38071 3893
rect 38286 3884 38292 3896
rect 38344 3884 38350 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 3142 3720 3148 3732
rect 2746 3692 3148 3720
rect 1765 3655 1823 3661
rect 1765 3621 1777 3655
rect 1811 3652 1823 3655
rect 2746 3652 2774 3692
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3252 3692 6500 3720
rect 3050 3652 3056 3664
rect 1811 3624 2774 3652
rect 3011 3624 3056 3652
rect 1811 3621 1823 3624
rect 1765 3615 1823 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 3252 3525 3280 3692
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3652 4951 3655
rect 5534 3652 5540 3664
rect 4939 3624 5540 3652
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 6472 3652 6500 3692
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 6972 3692 7389 3720
rect 6972 3680 6978 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 7484 3692 9904 3720
rect 7484 3652 7512 3692
rect 6472 3624 7512 3652
rect 7837 3655 7895 3661
rect 7837 3621 7849 3655
rect 7883 3652 7895 3655
rect 9876 3652 9904 3692
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 10284 3692 10333 3720
rect 10284 3680 10290 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10321 3683 10379 3689
rect 10428 3692 12572 3720
rect 10428 3652 10456 3692
rect 10781 3655 10839 3661
rect 10781 3652 10793 3655
rect 7883 3624 8064 3652
rect 9876 3624 10456 3652
rect 10520 3624 10793 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 3752 3556 5488 3584
rect 3752 3544 3758 3556
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2823 3488 3249 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 4890 3516 4896 3528
rect 4479 3488 4896 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 2424 3448 2452 3479
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 4982 3448 4988 3460
rect 2424 3420 4988 3448
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 5258 3380 5264 3392
rect 4295 3352 5264 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5460 3380 5488 3556
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 8036 3584 8064 3624
rect 8662 3584 8668 3596
rect 6604 3556 7954 3584
rect 8036 3556 8668 3584
rect 6604 3544 6610 3556
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 6362 3516 6368 3528
rect 5583 3488 6368 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 6362 3476 6368 3488
rect 6420 3516 6426 3528
rect 6822 3516 6828 3528
rect 6420 3488 6828 3516
rect 6420 3476 6426 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 5626 3408 5632 3460
rect 5684 3448 5690 3460
rect 5782 3451 5840 3457
rect 5782 3448 5794 3451
rect 5684 3420 5794 3448
rect 5684 3408 5690 3420
rect 5782 3417 5794 3420
rect 5828 3417 5840 3451
rect 7374 3448 7380 3460
rect 5782 3411 5840 3417
rect 6840 3420 7380 3448
rect 6840 3380 6868 3420
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7576 3448 7604 3479
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7926 3525 7954 3556
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 8846 3584 8852 3596
rect 8772 3556 8852 3584
rect 7883 3519 7954 3525
rect 7708 3488 7753 3516
rect 7708 3476 7714 3488
rect 7883 3485 7895 3519
rect 7929 3488 7954 3519
rect 8294 3516 8300 3528
rect 8036 3488 8300 3516
rect 7929 3485 7941 3488
rect 7883 3479 7941 3485
rect 8036 3448 8064 3488
rect 8294 3476 8300 3488
rect 8352 3516 8358 3528
rect 8772 3516 8800 3556
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10520 3584 10548 3624
rect 10781 3621 10793 3624
rect 10827 3621 10839 3655
rect 10781 3615 10839 3621
rect 11146 3584 11152 3596
rect 10284 3556 10548 3584
rect 10796 3556 11152 3584
rect 10284 3544 10290 3556
rect 8938 3516 8944 3528
rect 8352 3488 8800 3516
rect 8899 3488 8944 3516
rect 8352 3476 8358 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9197 3519 9255 3525
rect 9197 3516 9209 3519
rect 9088 3488 9209 3516
rect 9088 3476 9094 3488
rect 9197 3485 9209 3488
rect 9243 3485 9255 3519
rect 9197 3479 9255 3485
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 10796 3516 10824 3556
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 12544 3584 12572 3692
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12676 3692 12817 3720
rect 12676 3680 12682 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 14792 3692 15853 3720
rect 14792 3680 14798 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 15841 3683 15899 3689
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 18601 3723 18659 3729
rect 18601 3720 18613 3723
rect 16172 3692 18613 3720
rect 16172 3680 16178 3692
rect 18601 3689 18613 3692
rect 18647 3689 18659 3723
rect 21542 3720 21548 3732
rect 21503 3692 21548 3720
rect 18601 3683 18659 3689
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 22462 3720 22468 3732
rect 22112 3692 22468 3720
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 13265 3655 13323 3661
rect 13265 3652 13277 3655
rect 12768 3624 13277 3652
rect 12768 3612 12774 3624
rect 13265 3621 13277 3624
rect 13311 3621 13323 3655
rect 13265 3615 13323 3621
rect 13814 3584 13820 3596
rect 12544 3556 13820 3584
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 19242 3584 19248 3596
rect 19203 3556 19248 3584
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 22112 3593 22140 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23474 3720 23480 3732
rect 23435 3692 23480 3720
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 24765 3723 24823 3729
rect 24765 3689 24777 3723
rect 24811 3720 24823 3723
rect 26326 3720 26332 3732
rect 24811 3692 26332 3720
rect 24811 3689 24823 3692
rect 24765 3683 24823 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 26786 3720 26792 3732
rect 26747 3692 26792 3720
rect 26786 3680 26792 3692
rect 26844 3680 26850 3732
rect 28258 3720 28264 3732
rect 27639 3692 28264 3720
rect 22097 3587 22155 3593
rect 22097 3553 22109 3587
rect 22143 3553 22155 3587
rect 22097 3547 22155 3553
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 23256 3556 24409 3584
rect 23256 3544 23262 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 27639 3584 27667 3692
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 28997 3723 29055 3729
rect 28997 3689 29009 3723
rect 29043 3720 29055 3723
rect 29270 3720 29276 3732
rect 29043 3692 29276 3720
rect 29043 3689 29055 3692
rect 28997 3683 29055 3689
rect 29270 3680 29276 3692
rect 29328 3680 29334 3732
rect 29362 3680 29368 3732
rect 29420 3720 29426 3732
rect 29917 3723 29975 3729
rect 29420 3692 29776 3720
rect 29420 3680 29426 3692
rect 28810 3612 28816 3664
rect 28868 3652 28874 3664
rect 28868 3624 29592 3652
rect 28868 3612 28874 3624
rect 27639 3556 27752 3584
rect 24397 3547 24455 3553
rect 10962 3516 10968 3528
rect 9548 3488 10824 3516
rect 10923 3488 10968 3516
rect 9548 3476 9554 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 12158 3516 12164 3528
rect 11471 3488 12164 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 15194 3516 15200 3528
rect 14507 3488 15200 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 15194 3476 15200 3488
rect 15252 3516 15258 3528
rect 16390 3516 16396 3528
rect 15252 3488 16396 3516
rect 15252 3476 15258 3488
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 16649 3519 16707 3525
rect 16649 3516 16661 3519
rect 16540 3488 16661 3516
rect 16540 3476 16546 3488
rect 16649 3485 16661 3488
rect 16695 3485 16707 3519
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 16649 3479 16707 3485
rect 16776 3488 18245 3516
rect 16776 3460 16804 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 7576 3420 8064 3448
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 11146 3448 11152 3460
rect 8260 3420 11152 3448
rect 8260 3408 8266 3420
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11692 3451 11750 3457
rect 11692 3417 11704 3451
rect 11738 3448 11750 3451
rect 11974 3448 11980 3460
rect 11738 3420 11980 3448
rect 11738 3417 11750 3420
rect 11692 3411 11750 3417
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 14728 3451 14786 3457
rect 14728 3417 14740 3451
rect 14774 3448 14786 3451
rect 15746 3448 15752 3460
rect 14774 3420 15752 3448
rect 14774 3417 14786 3420
rect 14728 3411 14786 3417
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 16758 3408 16764 3460
rect 16816 3408 16822 3460
rect 17310 3408 17316 3460
rect 17368 3448 17374 3460
rect 18432 3448 18460 3479
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19501 3519 19559 3525
rect 19501 3516 19513 3519
rect 19392 3488 19513 3516
rect 19392 3476 19398 3488
rect 19501 3485 19513 3488
rect 19547 3485 19559 3519
rect 19501 3479 19559 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 21361 3519 21419 3525
rect 21361 3485 21373 3519
rect 21407 3516 21419 3519
rect 21726 3516 21732 3528
rect 21407 3488 21732 3516
rect 21407 3485 21419 3488
rect 21361 3479 21419 3485
rect 17368 3420 18460 3448
rect 17368 3408 17374 3420
rect 20990 3408 20996 3460
rect 21048 3448 21054 3460
rect 21284 3448 21312 3479
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 22364 3519 22422 3525
rect 22364 3485 22376 3519
rect 22410 3516 22422 3519
rect 22830 3516 22836 3528
rect 22410 3488 22836 3516
rect 22410 3485 22422 3488
rect 22364 3479 22422 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 24946 3516 24952 3528
rect 24627 3488 24952 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 25409 3519 25467 3525
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 27522 3516 27528 3528
rect 25455 3488 27528 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 27522 3476 27528 3488
rect 27580 3516 27586 3528
rect 27624 3519 27682 3525
rect 27624 3516 27636 3519
rect 27580 3488 27636 3516
rect 27580 3476 27586 3488
rect 27624 3485 27636 3488
rect 27670 3485 27682 3519
rect 27624 3479 27682 3485
rect 22186 3448 22192 3460
rect 21048 3420 22192 3448
rect 21048 3408 21054 3420
rect 22186 3408 22192 3420
rect 22244 3448 22250 3460
rect 25222 3448 25228 3460
rect 22244 3420 25228 3448
rect 22244 3408 22250 3420
rect 25222 3408 25228 3420
rect 25280 3408 25286 3460
rect 25676 3451 25734 3457
rect 25676 3417 25688 3451
rect 25722 3448 25734 3451
rect 27338 3448 27344 3460
rect 25722 3420 27344 3448
rect 25722 3417 25734 3420
rect 25676 3411 25734 3417
rect 27338 3408 27344 3420
rect 27396 3408 27402 3460
rect 27724 3448 27752 3556
rect 28718 3544 28724 3596
rect 28776 3584 28782 3596
rect 29270 3584 29276 3596
rect 28776 3556 29276 3584
rect 28776 3544 28782 3556
rect 29270 3544 29276 3556
rect 29328 3544 29334 3596
rect 29564 3593 29592 3624
rect 29549 3587 29607 3593
rect 29549 3553 29561 3587
rect 29595 3553 29607 3587
rect 29549 3547 29607 3553
rect 28166 3476 28172 3528
rect 28224 3516 28230 3528
rect 29748 3525 29776 3692
rect 29917 3689 29929 3723
rect 29963 3720 29975 3723
rect 33502 3720 33508 3732
rect 29963 3692 33508 3720
rect 29963 3689 29975 3692
rect 29917 3683 29975 3689
rect 33502 3680 33508 3692
rect 33560 3680 33566 3732
rect 33870 3680 33876 3732
rect 33928 3720 33934 3732
rect 34698 3720 34704 3732
rect 33928 3692 34704 3720
rect 33928 3680 33934 3692
rect 34698 3680 34704 3692
rect 34756 3680 34762 3732
rect 35897 3723 35955 3729
rect 35897 3689 35909 3723
rect 35943 3720 35955 3723
rect 36446 3720 36452 3732
rect 35943 3692 36452 3720
rect 35943 3689 35955 3692
rect 35897 3683 35955 3689
rect 36446 3680 36452 3692
rect 36504 3680 36510 3732
rect 34149 3655 34207 3661
rect 34149 3621 34161 3655
rect 34195 3652 34207 3655
rect 36630 3652 36636 3664
rect 34195 3624 36636 3652
rect 34195 3621 34207 3624
rect 34149 3615 34207 3621
rect 36630 3612 36636 3624
rect 36688 3612 36694 3664
rect 32306 3544 32312 3596
rect 32364 3584 32370 3596
rect 32950 3584 32956 3596
rect 32364 3556 32812 3584
rect 32911 3556 32956 3584
rect 32364 3544 32370 3556
rect 29733 3519 29791 3525
rect 28224 3488 29500 3516
rect 28224 3476 28230 3488
rect 27873 3451 27931 3457
rect 27873 3448 27885 3451
rect 27724 3420 27885 3448
rect 27873 3417 27885 3420
rect 27919 3417 27931 3451
rect 27873 3411 27931 3417
rect 27982 3408 27988 3460
rect 28040 3448 28046 3460
rect 29178 3448 29184 3460
rect 28040 3420 29184 3448
rect 28040 3408 28046 3420
rect 29178 3408 29184 3420
rect 29236 3408 29242 3460
rect 29472 3448 29500 3488
rect 29733 3485 29745 3519
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3516 30803 3519
rect 32214 3516 32220 3528
rect 30791 3488 32220 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 32214 3476 32220 3488
rect 32272 3516 32278 3528
rect 32398 3516 32404 3528
rect 32272 3488 32404 3516
rect 32272 3476 32278 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 32784 3525 32812 3556
rect 32950 3544 32956 3556
rect 33008 3544 33014 3596
rect 33042 3544 33048 3596
rect 33100 3584 33106 3596
rect 33781 3587 33839 3593
rect 33100 3556 33272 3584
rect 33100 3544 33106 3556
rect 32585 3519 32643 3525
rect 32585 3485 32597 3519
rect 32631 3485 32643 3519
rect 32585 3479 32643 3485
rect 32769 3519 32827 3525
rect 32769 3485 32781 3519
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 32861 3519 32919 3525
rect 32861 3485 32873 3519
rect 32907 3485 32919 3519
rect 33134 3516 33140 3528
rect 33095 3488 33140 3516
rect 32861 3479 32919 3485
rect 30650 3448 30656 3460
rect 29472 3420 30656 3448
rect 30650 3408 30656 3420
rect 30708 3408 30714 3460
rect 31012 3451 31070 3457
rect 31012 3417 31024 3451
rect 31058 3448 31070 3451
rect 31386 3448 31392 3460
rect 31058 3420 31392 3448
rect 31058 3417 31070 3420
rect 31012 3411 31070 3417
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 31478 3408 31484 3460
rect 31536 3448 31542 3460
rect 31536 3420 31616 3448
rect 31536 3408 31542 3420
rect 5460 3352 6868 3380
rect 6917 3383 6975 3389
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 7650 3380 7656 3392
rect 6963 3352 7656 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 10502 3380 10508 3392
rect 7892 3352 10508 3380
rect 7892 3340 7898 3352
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 17770 3380 17776 3392
rect 17731 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 20622 3380 20628 3392
rect 20583 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 30834 3380 30840 3392
rect 24912 3352 30840 3380
rect 24912 3340 24918 3352
rect 30834 3340 30840 3352
rect 30892 3340 30898 3392
rect 31588 3380 31616 3420
rect 32306 3408 32312 3460
rect 32364 3448 32370 3460
rect 32600 3448 32628 3479
rect 32364 3420 32628 3448
rect 32876 3448 32904 3479
rect 33134 3476 33140 3488
rect 33192 3476 33198 3528
rect 33244 3516 33272 3556
rect 33781 3553 33793 3587
rect 33827 3584 33839 3587
rect 34701 3587 34759 3593
rect 34701 3584 34713 3587
rect 33827 3556 34713 3584
rect 33827 3553 33839 3556
rect 33781 3547 33839 3553
rect 34701 3553 34713 3556
rect 34747 3584 34759 3587
rect 34974 3584 34980 3596
rect 34747 3556 34980 3584
rect 34747 3553 34759 3556
rect 34701 3547 34759 3553
rect 34974 3544 34980 3556
rect 35032 3584 35038 3596
rect 35529 3587 35587 3593
rect 35529 3584 35541 3587
rect 35032 3556 35541 3584
rect 35032 3544 35038 3556
rect 35529 3553 35541 3556
rect 35575 3584 35587 3587
rect 35618 3584 35624 3596
rect 35575 3556 35624 3584
rect 35575 3553 35587 3556
rect 35529 3547 35587 3553
rect 35618 3544 35624 3556
rect 35676 3544 35682 3596
rect 33965 3519 34023 3525
rect 33965 3516 33977 3519
rect 33244 3488 33977 3516
rect 33965 3485 33977 3488
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34848 3488 34897 3516
rect 34848 3476 34854 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 35710 3516 35716 3528
rect 35671 3488 35716 3516
rect 34885 3479 34943 3485
rect 35710 3476 35716 3488
rect 35768 3476 35774 3528
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 36357 3519 36415 3525
rect 36357 3516 36369 3519
rect 36228 3488 36369 3516
rect 36228 3476 36234 3488
rect 36357 3485 36369 3488
rect 36403 3485 36415 3519
rect 36357 3479 36415 3485
rect 37645 3519 37703 3525
rect 37645 3485 37657 3519
rect 37691 3485 37703 3519
rect 37645 3479 37703 3485
rect 33226 3448 33232 3460
rect 32876 3420 33232 3448
rect 32364 3408 32370 3420
rect 32125 3383 32183 3389
rect 32125 3380 32137 3383
rect 31588 3352 32137 3380
rect 32125 3349 32137 3352
rect 32171 3349 32183 3383
rect 32125 3343 32183 3349
rect 32582 3340 32588 3392
rect 32640 3380 32646 3392
rect 32876 3380 32904 3420
rect 33226 3408 33232 3420
rect 33284 3408 33290 3460
rect 33321 3451 33379 3457
rect 33321 3417 33333 3451
rect 33367 3448 33379 3451
rect 37660 3448 37688 3479
rect 33367 3420 37688 3448
rect 33367 3417 33379 3420
rect 33321 3411 33379 3417
rect 32640 3352 32904 3380
rect 32640 3340 32646 3352
rect 34514 3340 34520 3392
rect 34572 3380 34578 3392
rect 34790 3380 34796 3392
rect 34572 3352 34796 3380
rect 34572 3340 34578 3352
rect 34790 3340 34796 3352
rect 34848 3340 34854 3392
rect 35069 3383 35127 3389
rect 35069 3349 35081 3383
rect 35115 3380 35127 3383
rect 35802 3380 35808 3392
rect 35115 3352 35808 3380
rect 35115 3349 35127 3352
rect 35069 3343 35127 3349
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 36078 3340 36084 3392
rect 36136 3380 36142 3392
rect 36541 3383 36599 3389
rect 36541 3380 36553 3383
rect 36136 3352 36553 3380
rect 36136 3340 36142 3352
rect 36541 3349 36553 3352
rect 36587 3349 36599 3383
rect 36541 3343 36599 3349
rect 37550 3340 37556 3392
rect 37608 3380 37614 3392
rect 37829 3383 37887 3389
rect 37829 3380 37841 3383
rect 37608 3352 37841 3380
rect 37608 3340 37614 3352
rect 37829 3349 37841 3352
rect 37875 3349 37887 3383
rect 37829 3343 37887 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2067 3179 2125 3185
rect 2067 3145 2079 3179
rect 2113 3176 2125 3179
rect 2682 3176 2688 3188
rect 2113 3148 2688 3176
rect 2113 3145 2125 3148
rect 2067 3139 2125 3145
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3234 3176 3240 3188
rect 3099 3148 3240 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4387 3148 5580 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 1854 3108 1860 3120
rect 1815 3080 1860 3108
rect 1854 3068 1860 3080
rect 1912 3068 1918 3120
rect 5442 3108 5448 3120
rect 4540 3080 5448 3108
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4430 3040 4436 3052
rect 3927 3012 4436 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3252 2972 3280 3003
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4540 3049 4568 3080
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 5552 3108 5580 3148
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 5684 3148 5729 3176
rect 5684 3136 5690 3148
rect 6546 3136 6552 3188
rect 6604 3136 6610 3188
rect 7834 3136 7840 3188
rect 7892 3136 7898 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 10318 3176 10324 3188
rect 8076 3148 10324 3176
rect 8076 3136 8082 3148
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 10686 3136 10692 3188
rect 10744 3176 10750 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10744 3148 10977 3176
rect 10744 3136 10750 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 13630 3176 13636 3188
rect 11204 3148 13636 3176
rect 11204 3136 11210 3148
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14568 3148 15056 3176
rect 6564 3108 6592 3136
rect 6638 3117 6644 3120
rect 5552 3080 6592 3108
rect 6632 3071 6644 3117
rect 6696 3108 6702 3120
rect 7852 3108 7880 3136
rect 6696 3080 6732 3108
rect 7852 3080 8616 3108
rect 6638 3068 6644 3071
rect 6696 3068 6702 3080
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5534 3040 5540 3052
rect 5215 3012 5540 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7190 3040 7196 3052
rect 6472 3012 7196 3040
rect 4614 2972 4620 2984
rect 3252 2944 4620 2972
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 6472 2972 6500 3012
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8588 3049 8616 3080
rect 8938 3068 8944 3120
rect 8996 3108 9002 3120
rect 12158 3108 12164 3120
rect 8996 3080 12164 3108
rect 8996 3068 9002 3080
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8352 3012 8401 3040
rect 8352 3000 8358 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8541 3043 8616 3049
rect 8541 3009 8553 3043
rect 8587 3012 8616 3043
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8587 3009 8599 3012
rect 8541 3003 8599 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9600 3049 9628 3080
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9674 3000 9680 3052
rect 9732 3000 9738 3052
rect 9852 3043 9910 3049
rect 9852 3009 9864 3043
rect 9898 3040 9910 3043
rect 10226 3040 10232 3052
rect 9898 3012 10232 3040
rect 9898 3009 9910 3012
rect 9852 3003 9910 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11808 3049 11836 3080
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 13906 3108 13912 3120
rect 13867 3080 13912 3108
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 12066 3049 12072 3052
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 12060 3003 12072 3049
rect 12124 3040 12130 3052
rect 12124 3012 12160 3040
rect 12066 3000 12072 3003
rect 12124 3000 12130 3012
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 13228 3012 13645 3040
rect 13228 3000 13234 3012
rect 13633 3009 13645 3012
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13780 3012 13829 3040
rect 13780 3000 13786 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3040 14059 3043
rect 14568 3040 14596 3148
rect 14918 3108 14924 3120
rect 14879 3080 14924 3108
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 14047 3012 14596 3040
rect 14645 3043 14703 3049
rect 14047 3009 14059 3012
rect 14001 3003 14059 3009
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 9692 2972 9720 3000
rect 5000 2944 6500 2972
rect 8128 2944 9720 2972
rect 13832 2972 13860 3003
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15028 3049 15056 3148
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 16724 3148 18061 3176
rect 16724 3136 16730 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 19981 3179 20039 3185
rect 19981 3145 19993 3179
rect 20027 3176 20039 3179
rect 20438 3176 20444 3188
rect 20027 3148 20444 3176
rect 20027 3145 20039 3148
rect 19981 3139 20039 3145
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 20956 3148 21281 3176
rect 20956 3136 20962 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 21269 3139 21327 3145
rect 22051 3179 22109 3185
rect 22051 3145 22063 3179
rect 22097 3145 22109 3179
rect 22051 3139 22109 3145
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 16758 3108 16764 3120
rect 15764 3080 16764 3108
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15286 3040 15292 3052
rect 15059 3012 15292 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 14844 2972 14872 3003
rect 15286 3000 15292 3012
rect 15344 3000 15350 3052
rect 15764 3049 15792 3080
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 15102 2972 15108 2984
rect 13832 2944 15108 2972
rect 2222 2904 2228 2916
rect 2183 2876 2228 2904
rect 2222 2864 2228 2876
rect 2280 2864 2286 2916
rect 5000 2913 5028 2944
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2873 5043 2907
rect 4985 2867 5043 2873
rect 7650 2864 7656 2916
rect 7708 2904 7714 2916
rect 7745 2907 7803 2913
rect 7745 2904 7757 2907
rect 7708 2876 7757 2904
rect 7708 2864 7714 2876
rect 7745 2873 7757 2876
rect 7791 2873 7803 2907
rect 8128 2904 8156 2944
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15856 2972 15884 3003
rect 15212 2944 15884 2972
rect 8662 2904 8668 2916
rect 7745 2867 7803 2873
rect 7843 2876 8156 2904
rect 8575 2876 8668 2904
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 4062 2836 4068 2848
rect 3743 2808 4068 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 7843 2836 7871 2876
rect 8662 2864 8668 2876
rect 8720 2904 8726 2916
rect 9582 2904 9588 2916
rect 8720 2876 9588 2904
rect 8720 2864 8726 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 14090 2904 14096 2916
rect 13096 2876 14096 2904
rect 5132 2808 7871 2836
rect 5132 2796 5138 2808
rect 7926 2796 7932 2848
rect 7984 2836 7990 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7984 2808 8217 2836
rect 7984 2796 7990 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 10594 2836 10600 2848
rect 8996 2808 10600 2836
rect 8996 2796 9002 2808
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 13096 2836 13124 2876
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 15212 2913 15240 2944
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2873 15255 2907
rect 15948 2904 15976 3080
rect 16758 3068 16764 3080
rect 16816 3068 16822 3120
rect 16936 3111 16994 3117
rect 16936 3077 16948 3111
rect 16982 3108 16994 3111
rect 17218 3108 17224 3120
rect 16982 3080 17224 3108
rect 16982 3077 16994 3080
rect 16936 3071 16994 3077
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 22066 3108 22094 3139
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 25774 3136 25780 3188
rect 25832 3176 25838 3188
rect 26329 3179 26387 3185
rect 26329 3176 26341 3179
rect 25832 3148 26341 3176
rect 25832 3136 25838 3148
rect 26329 3145 26341 3148
rect 26375 3145 26387 3179
rect 26329 3139 26387 3145
rect 27798 3136 27804 3188
rect 27856 3176 27862 3188
rect 30466 3176 30472 3188
rect 27856 3148 30472 3176
rect 27856 3136 27862 3148
rect 30466 3136 30472 3148
rect 30524 3136 30530 3188
rect 30668 3148 32444 3176
rect 28166 3108 28172 3120
rect 19116 3080 22094 3108
rect 23032 3080 24900 3108
rect 19116 3068 19122 3080
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16448 3012 16681 3040
rect 16448 3000 16454 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 19150 3040 19156 3052
rect 18555 3012 19156 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 19150 3000 19156 3012
rect 19208 3000 19214 3052
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20622 3040 20628 3052
rect 19751 3012 20628 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20990 3040 20996 3052
rect 20951 3012 20996 3040
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3040 21143 3043
rect 22370 3040 22376 3052
rect 21131 3012 22376 3040
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20346 2972 20352 2984
rect 20027 2944 20352 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 21818 2972 21824 2984
rect 21779 2944 21824 2972
rect 21818 2932 21824 2944
rect 21876 2972 21882 2984
rect 23032 2972 23060 3080
rect 24872 3052 24900 3080
rect 25056 3080 28172 3108
rect 23198 3040 23204 3052
rect 23159 3012 23204 3040
rect 23198 3000 23204 3012
rect 23256 3000 23262 3052
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 24121 3043 24179 3049
rect 23348 3012 23393 3040
rect 23348 3000 23354 3012
rect 24121 3009 24133 3043
rect 24167 3040 24179 3043
rect 24578 3040 24584 3052
rect 24167 3012 24584 3040
rect 24167 3009 24179 3012
rect 24121 3003 24179 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 24854 3040 24860 3052
rect 24815 3012 24860 3040
rect 24854 3000 24860 3012
rect 24912 3000 24918 3052
rect 21876 2944 23060 2972
rect 21876 2932 21882 2944
rect 15197 2867 15255 2873
rect 15304 2876 15976 2904
rect 19797 2907 19855 2913
rect 12032 2808 13124 2836
rect 12032 2796 12038 2808
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 13228 2808 13273 2836
rect 13228 2796 13234 2808
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 14274 2836 14280 2848
rect 13872 2808 14280 2836
rect 13872 2796 13878 2808
rect 14274 2796 14280 2808
rect 14332 2836 14338 2848
rect 15304 2836 15332 2876
rect 19797 2873 19809 2907
rect 19843 2904 19855 2907
rect 25056 2904 25084 3080
rect 28166 3068 28172 3080
rect 28224 3068 28230 3120
rect 28445 3111 28503 3117
rect 28445 3077 28457 3111
rect 28491 3108 28503 3111
rect 29273 3111 29331 3117
rect 28491 3080 29224 3108
rect 28491 3077 28503 3080
rect 28445 3071 28503 3077
rect 25133 3043 25191 3049
rect 25133 3009 25145 3043
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25148 2972 25176 3003
rect 25958 3000 25964 3052
rect 26016 3040 26022 3052
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 26016 3012 26249 3040
rect 26016 3000 26022 3012
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 26237 3003 26295 3009
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 27706 3040 27712 3052
rect 27540 3012 27712 3040
rect 26510 2972 26516 2984
rect 25148 2944 26516 2972
rect 26510 2932 26516 2944
rect 26568 2932 26574 2984
rect 27249 2975 27307 2981
rect 27249 2941 27261 2975
rect 27295 2972 27307 2975
rect 27540 2972 27568 3012
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 27890 3000 27896 3052
rect 27948 3040 27954 3052
rect 28261 3043 28319 3049
rect 28261 3040 28273 3043
rect 27948 3012 28273 3040
rect 27948 3000 27954 3012
rect 28261 3009 28273 3012
rect 28307 3009 28319 3043
rect 28261 3003 28319 3009
rect 28350 3000 28356 3052
rect 28408 3040 28414 3052
rect 29089 3043 29147 3049
rect 29089 3040 29101 3043
rect 28408 3012 29101 3040
rect 28408 3000 28414 3012
rect 29089 3009 29101 3012
rect 29135 3009 29147 3043
rect 29089 3003 29147 3009
rect 27295 2944 27568 2972
rect 27617 2975 27675 2981
rect 27295 2941 27307 2944
rect 27249 2935 27307 2941
rect 27617 2941 27629 2975
rect 27663 2972 27675 2975
rect 27982 2972 27988 2984
rect 27663 2944 27988 2972
rect 27663 2941 27675 2944
rect 27617 2935 27675 2941
rect 27982 2932 27988 2944
rect 28040 2932 28046 2984
rect 28077 2975 28135 2981
rect 28077 2941 28089 2975
rect 28123 2972 28135 2975
rect 28810 2972 28816 2984
rect 28123 2944 28816 2972
rect 28123 2941 28135 2944
rect 28077 2935 28135 2941
rect 28810 2932 28816 2944
rect 28868 2972 28874 2984
rect 28905 2975 28963 2981
rect 28905 2972 28917 2975
rect 28868 2944 28917 2972
rect 28868 2932 28874 2944
rect 28905 2941 28917 2944
rect 28951 2941 28963 2975
rect 29196 2972 29224 3080
rect 29273 3077 29285 3111
rect 29319 3108 29331 3111
rect 30668 3108 30696 3148
rect 29319 3080 30696 3108
rect 32416 3108 32444 3148
rect 32490 3136 32496 3188
rect 32548 3176 32554 3188
rect 34514 3176 34520 3188
rect 32548 3148 34520 3176
rect 32548 3136 32554 3148
rect 34514 3136 34520 3148
rect 34572 3136 34578 3188
rect 36354 3176 36360 3188
rect 34624 3148 36360 3176
rect 32416 3080 34468 3108
rect 29319 3077 29331 3080
rect 29273 3071 29331 3077
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 30834 3040 30840 3052
rect 30795 3012 30840 3040
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 30926 3000 30932 3052
rect 30984 3040 30990 3052
rect 31021 3043 31079 3049
rect 31021 3040 31033 3043
rect 30984 3012 31033 3040
rect 30984 3000 30990 3012
rect 31021 3009 31033 3012
rect 31067 3009 31079 3043
rect 31021 3003 31079 3009
rect 31110 3000 31116 3052
rect 31168 3040 31174 3052
rect 31168 3012 31213 3040
rect 31168 3000 31174 3012
rect 31294 3000 31300 3052
rect 31352 3040 31358 3052
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 31352 3012 31401 3040
rect 31352 3000 31358 3012
rect 31389 3009 31401 3012
rect 31435 3009 31447 3043
rect 32398 3040 32404 3052
rect 32359 3012 32404 3040
rect 31389 3003 31447 3009
rect 32398 3000 32404 3012
rect 32456 3000 32462 3052
rect 32674 3049 32680 3052
rect 32668 3040 32680 3049
rect 32635 3012 32680 3040
rect 32668 3003 32680 3012
rect 32674 3000 32680 3003
rect 32732 3000 32738 3052
rect 34440 3049 34468 3080
rect 34425 3043 34483 3049
rect 34425 3009 34437 3043
rect 34471 3009 34483 3043
rect 34425 3003 34483 3009
rect 29822 2972 29828 2984
rect 29196 2944 29828 2972
rect 28905 2935 28963 2941
rect 29822 2932 29828 2944
rect 29880 2932 29886 2984
rect 31202 2972 31208 2984
rect 31115 2944 31208 2972
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 33778 2932 33784 2984
rect 33836 2972 33842 2984
rect 34624 2972 34652 3148
rect 36354 3136 36360 3148
rect 36412 3136 36418 3188
rect 34790 3068 34796 3120
rect 34848 3108 34854 3120
rect 34848 3080 35112 3108
rect 34848 3068 34854 3080
rect 34974 3040 34980 3052
rect 34935 3012 34980 3040
rect 34974 3000 34980 3012
rect 35032 3000 35038 3052
rect 35084 3049 35112 3080
rect 35802 3068 35808 3120
rect 35860 3108 35866 3120
rect 35860 3080 36768 3108
rect 35860 3068 35866 3080
rect 35069 3043 35127 3049
rect 35069 3009 35081 3043
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35253 3043 35311 3049
rect 35253 3009 35265 3043
rect 35299 3040 35311 3043
rect 35897 3043 35955 3049
rect 35299 3012 35848 3040
rect 35299 3009 35311 3012
rect 35253 3003 35311 3009
rect 33836 2944 34652 2972
rect 33836 2932 33842 2944
rect 35434 2932 35440 2984
rect 35492 2972 35498 2984
rect 35713 2975 35771 2981
rect 35713 2972 35725 2975
rect 35492 2944 35725 2972
rect 35492 2932 35498 2944
rect 35713 2941 35725 2944
rect 35759 2941 35771 2975
rect 35820 2972 35848 3012
rect 35897 3009 35909 3043
rect 35943 3040 35955 3043
rect 35986 3040 35992 3052
rect 35943 3012 35992 3040
rect 35943 3009 35955 3012
rect 35897 3003 35955 3009
rect 35986 3000 35992 3012
rect 36044 3000 36050 3052
rect 36081 3043 36139 3049
rect 36081 3009 36093 3043
rect 36127 3040 36139 3043
rect 36630 3040 36636 3052
rect 36127 3012 36636 3040
rect 36127 3009 36139 3012
rect 36081 3003 36139 3009
rect 36630 3000 36636 3012
rect 36688 3000 36694 3052
rect 36740 3049 36768 3080
rect 36725 3043 36783 3049
rect 36725 3009 36737 3043
rect 36771 3009 36783 3043
rect 37274 3040 37280 3052
rect 37235 3012 37280 3040
rect 36725 3003 36783 3009
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 36538 2972 36544 2984
rect 35820 2944 36544 2972
rect 35713 2935 35771 2941
rect 36538 2932 36544 2944
rect 36596 2932 36602 2984
rect 37458 2932 37464 2984
rect 37516 2932 37522 2984
rect 19843 2876 25084 2904
rect 19843 2873 19855 2876
rect 19797 2867 19855 2873
rect 27062 2864 27068 2916
rect 27120 2904 27126 2916
rect 28994 2904 29000 2916
rect 27120 2876 29000 2904
rect 27120 2864 27126 2876
rect 28994 2864 29000 2876
rect 29052 2864 29058 2916
rect 29917 2907 29975 2913
rect 29917 2904 29929 2907
rect 29104 2876 29929 2904
rect 16022 2836 16028 2848
rect 14332 2808 15332 2836
rect 15983 2808 16028 2836
rect 14332 2796 14338 2808
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18693 2839 18751 2845
rect 18693 2836 18705 2839
rect 18196 2808 18705 2836
rect 18196 2796 18202 2808
rect 18693 2805 18705 2808
rect 18739 2805 18751 2839
rect 18693 2799 18751 2805
rect 21818 2796 21824 2848
rect 21876 2836 21882 2848
rect 23106 2836 23112 2848
rect 21876 2808 23112 2836
rect 21876 2796 21882 2808
rect 23106 2796 23112 2808
rect 23164 2796 23170 2848
rect 24305 2839 24363 2845
rect 24305 2805 24317 2839
rect 24351 2836 24363 2839
rect 24854 2836 24860 2848
rect 24351 2808 24860 2836
rect 24351 2805 24363 2808
rect 24305 2799 24363 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25222 2796 25228 2848
rect 25280 2836 25286 2848
rect 28166 2836 28172 2848
rect 25280 2808 28172 2836
rect 25280 2796 25286 2808
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 28534 2796 28540 2848
rect 28592 2836 28598 2848
rect 29104 2836 29132 2876
rect 29917 2873 29929 2876
rect 29963 2873 29975 2907
rect 29917 2867 29975 2873
rect 28592 2808 29132 2836
rect 28592 2796 28598 2808
rect 29270 2796 29276 2848
rect 29328 2836 29334 2848
rect 31220 2836 31248 2932
rect 33410 2864 33416 2916
rect 33468 2904 33474 2916
rect 34241 2907 34299 2913
rect 34241 2904 34253 2907
rect 33468 2876 34253 2904
rect 33468 2864 33474 2876
rect 34241 2873 34253 2876
rect 34287 2873 34299 2907
rect 34241 2867 34299 2873
rect 34790 2864 34796 2916
rect 34848 2904 34854 2916
rect 37476 2904 37504 2932
rect 34848 2876 37504 2904
rect 34848 2864 34854 2876
rect 29328 2808 31248 2836
rect 31573 2839 31631 2845
rect 29328 2796 29334 2808
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 32766 2836 32772 2848
rect 31619 2808 32772 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 32766 2796 32772 2808
rect 32824 2796 32830 2848
rect 33134 2796 33140 2848
rect 33192 2836 33198 2848
rect 33781 2839 33839 2845
rect 33781 2836 33793 2839
rect 33192 2808 33793 2836
rect 33192 2796 33198 2808
rect 33781 2805 33793 2808
rect 33827 2805 33839 2839
rect 33781 2799 33839 2805
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36541 2839 36599 2845
rect 36541 2836 36553 2839
rect 36228 2808 36553 2836
rect 36228 2796 36234 2808
rect 36541 2805 36553 2808
rect 36587 2805 36599 2839
rect 36541 2799 36599 2805
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36872 2808 37473 2836
rect 36872 2796 36878 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6638 2632 6644 2644
rect 6411 2604 6644 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 8110 2632 8116 2644
rect 7432 2604 7604 2632
rect 8071 2604 8116 2632
rect 7432 2592 7438 2604
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2130 2564 2136 2576
rect 2087 2536 2136 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 2130 2524 2136 2536
rect 2188 2524 2194 2576
rect 4706 2524 4712 2576
rect 4764 2524 4770 2576
rect 5166 2524 5172 2576
rect 5224 2564 5230 2576
rect 7466 2564 7472 2576
rect 5224 2536 7472 2564
rect 5224 2524 5230 2536
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 4724 2496 4752 2524
rect 6914 2496 6920 2508
rect 4724 2468 6920 2496
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7576 2496 7604 2604
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9306 2632 9312 2644
rect 9267 2604 9312 2632
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10962 2632 10968 2644
rect 10459 2604 10968 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 15838 2632 15844 2644
rect 15799 2604 15844 2632
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 18690 2632 18696 2644
rect 17083 2604 18696 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 22186 2592 22192 2644
rect 22244 2632 22250 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 22244 2604 22385 2632
rect 22244 2592 22250 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 22373 2595 22431 2601
rect 26053 2635 26111 2641
rect 26053 2601 26065 2635
rect 26099 2632 26111 2635
rect 28074 2632 28080 2644
rect 26099 2604 28080 2632
rect 26099 2601 26111 2604
rect 26053 2595 26111 2601
rect 28074 2592 28080 2604
rect 28132 2592 28138 2644
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28813 2635 28871 2641
rect 28813 2632 28825 2635
rect 28408 2604 28825 2632
rect 28408 2592 28414 2604
rect 28813 2601 28825 2604
rect 28859 2601 28871 2635
rect 28813 2595 28871 2601
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 17310 2564 17316 2576
rect 15427 2536 17316 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 17310 2524 17316 2536
rect 17368 2524 17374 2576
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 17460 2536 18429 2564
rect 17460 2524 17466 2536
rect 18417 2533 18429 2536
rect 18463 2533 18475 2567
rect 18417 2527 18475 2533
rect 21082 2524 21088 2576
rect 21140 2564 21146 2576
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 21140 2536 23121 2564
rect 21140 2524 21146 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 23109 2527 23167 2533
rect 25590 2524 25596 2576
rect 25648 2564 25654 2576
rect 27157 2567 27215 2573
rect 27157 2564 27169 2567
rect 25648 2536 27169 2564
rect 25648 2524 25654 2536
rect 27157 2533 27169 2536
rect 27203 2533 27215 2567
rect 28828 2564 28856 2595
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 29052 2604 29745 2632
rect 29052 2592 29058 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 30466 2632 30472 2644
rect 30427 2604 30472 2632
rect 29733 2595 29791 2601
rect 30466 2592 30472 2604
rect 30524 2592 30530 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 31588 2604 32321 2632
rect 29270 2564 29276 2576
rect 28828 2536 29276 2564
rect 27157 2527 27215 2533
rect 29270 2524 29276 2536
rect 29328 2524 29334 2576
rect 29362 2524 29368 2576
rect 29420 2564 29426 2576
rect 31205 2567 31263 2573
rect 31205 2564 31217 2567
rect 29420 2536 31217 2564
rect 29420 2524 29426 2536
rect 31205 2533 31217 2536
rect 31251 2533 31263 2567
rect 31205 2527 31263 2533
rect 13998 2496 14004 2508
rect 7576 2468 11100 2496
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 3936 2400 4721 2428
rect 3936 2388 3942 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 6595 2400 7389 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 624 2332 1869 2360
rect 624 2320 630 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 4246 2320 4252 2372
rect 4304 2360 4310 2372
rect 5368 2360 5396 2391
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 8076 2400 8309 2428
rect 8076 2388 8082 2400
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 9398 2428 9404 2440
rect 8987 2400 9404 2428
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10410 2428 10416 2440
rect 10091 2400 10416 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10962 2388 10968 2440
rect 11020 2388 11026 2440
rect 4304 2332 5396 2360
rect 7009 2363 7067 2369
rect 4304 2320 4310 2332
rect 7009 2329 7021 2363
rect 7055 2329 7067 2363
rect 7009 2323 7067 2329
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3200 2264 3985 2292
rect 3200 2252 3206 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 3973 2255 4031 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 7024 2292 7052 2323
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7193 2363 7251 2369
rect 7193 2360 7205 2363
rect 7156 2332 7205 2360
rect 7156 2320 7162 2332
rect 7193 2329 7205 2332
rect 7239 2360 7251 2363
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 7239 2332 9137 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 9125 2329 9137 2332
rect 9171 2360 9183 2363
rect 10229 2363 10287 2369
rect 10229 2360 10241 2363
rect 9171 2332 10241 2360
rect 9171 2329 9183 2332
rect 9125 2323 9183 2329
rect 10229 2329 10241 2332
rect 10275 2360 10287 2363
rect 10980 2360 11008 2388
rect 10275 2332 11008 2360
rect 10275 2329 10287 2332
rect 10229 2323 10287 2329
rect 7926 2292 7932 2304
rect 7024 2264 7932 2292
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 11072 2292 11100 2468
rect 12406 2468 14004 2496
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12406 2428 12434 2468
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 17770 2496 17776 2508
rect 14844 2468 17776 2496
rect 14844 2440 14872 2468
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 25498 2456 25504 2508
rect 25556 2496 25562 2508
rect 28442 2496 28448 2508
rect 25556 2468 25912 2496
rect 25556 2456 25562 2468
rect 12299 2400 12434 2428
rect 12713 2431 12771 2437
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 12713 2391 12771 2397
rect 12728 2360 12756 2391
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13127 2400 14289 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14826 2428 14832 2440
rect 14787 2400 14832 2428
rect 14277 2391 14335 2397
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 15010 2428 15016 2440
rect 14971 2400 15016 2428
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15286 2428 15292 2440
rect 15243 2400 15292 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 17954 2428 17960 2440
rect 17543 2400 17960 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18230 2428 18236 2440
rect 18191 2400 18236 2428
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19426 2428 19432 2440
rect 19291 2400 19432 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19978 2428 19984 2440
rect 19939 2400 19984 2428
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20714 2428 20720 2440
rect 20675 2400 20720 2428
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 22922 2428 22928 2440
rect 22883 2400 22928 2428
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 25038 2428 25044 2440
rect 24443 2400 25044 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25884 2437 25912 2468
rect 26988 2468 28448 2496
rect 26988 2437 27016 2468
rect 28442 2456 28448 2468
rect 28500 2456 28506 2508
rect 29638 2496 29644 2508
rect 28736 2468 29644 2496
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25188 2400 25697 2428
rect 25188 2388 25194 2400
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2428 27767 2431
rect 28736 2428 28764 2468
rect 29638 2456 29644 2468
rect 29696 2456 29702 2508
rect 30098 2456 30104 2508
rect 30156 2496 30162 2508
rect 31588 2496 31616 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 34514 2592 34520 2644
rect 34572 2632 34578 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34572 2604 34897 2632
rect 34572 2592 34578 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 36354 2632 36360 2644
rect 36315 2604 36360 2632
rect 34885 2595 34943 2601
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 37458 2632 37464 2644
rect 37419 2604 37464 2632
rect 37458 2592 37464 2604
rect 37516 2592 37522 2644
rect 31662 2524 31668 2576
rect 31720 2564 31726 2576
rect 33781 2567 33839 2573
rect 33781 2564 33793 2567
rect 31720 2536 33793 2564
rect 31720 2524 31726 2536
rect 33781 2533 33793 2536
rect 33827 2533 33839 2567
rect 33781 2527 33839 2533
rect 30156 2468 31616 2496
rect 30156 2456 30162 2468
rect 32766 2456 32772 2508
rect 32824 2496 32830 2508
rect 32824 2468 33640 2496
rect 32824 2456 32830 2468
rect 29546 2428 29552 2440
rect 27755 2400 28764 2428
rect 29507 2400 29552 2428
rect 27755 2397 27767 2400
rect 27709 2391 27767 2397
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 30190 2388 30196 2440
rect 30248 2428 30254 2440
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 30248 2400 30297 2428
rect 30248 2388 30254 2400
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 31018 2428 31024 2440
rect 30979 2400 31024 2428
rect 30285 2391 30343 2397
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31628 2400 32137 2428
rect 31628 2388 31634 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33410 2428 33416 2440
rect 32907 2400 33416 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33410 2388 33416 2400
rect 33468 2388 33474 2440
rect 33612 2437 33640 2468
rect 34606 2456 34612 2508
rect 34664 2496 34670 2508
rect 34664 2468 35480 2496
rect 34664 2456 34670 2468
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 34698 2428 34704 2440
rect 34659 2400 34704 2428
rect 33597 2391 33655 2397
rect 34698 2388 34704 2400
rect 34756 2388 34762 2440
rect 35452 2437 35480 2468
rect 35437 2431 35495 2437
rect 35437 2397 35449 2431
rect 35483 2397 35495 2431
rect 36170 2428 36176 2440
rect 36131 2400 36176 2428
rect 35437 2391 35495 2397
rect 36170 2388 36176 2400
rect 36228 2388 36234 2440
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2428 37335 2431
rect 37366 2428 37372 2440
rect 37323 2400 37372 2428
rect 37323 2397 37335 2400
rect 37277 2391 37335 2397
rect 37366 2388 37372 2400
rect 37424 2388 37430 2440
rect 13814 2360 13820 2372
rect 12728 2332 13820 2360
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 15105 2363 15163 2369
rect 15105 2329 15117 2363
rect 15151 2329 15163 2363
rect 15105 2323 15163 2329
rect 15120 2292 15148 2323
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 22281 2363 22339 2369
rect 16632 2332 17724 2360
rect 16632 2320 16638 2332
rect 17696 2301 17724 2332
rect 22281 2329 22293 2363
rect 22327 2360 22339 2363
rect 22646 2360 22652 2372
rect 22327 2332 22652 2360
rect 22327 2329 22339 2332
rect 22281 2323 22339 2329
rect 22646 2320 22652 2332
rect 22704 2320 22710 2372
rect 28626 2320 28632 2372
rect 28684 2360 28690 2372
rect 28721 2363 28779 2369
rect 28721 2360 28733 2363
rect 28684 2332 28733 2360
rect 28684 2320 28690 2332
rect 28721 2329 28733 2332
rect 28767 2329 28779 2363
rect 28721 2323 28779 2329
rect 11072 2264 15148 2292
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 18874 2252 18880 2304
rect 18932 2292 18938 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18932 2264 19441 2292
rect 18932 2252 18938 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20036 2264 20177 2292
rect 20036 2252 20042 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20346 2252 20352 2304
rect 20404 2292 20410 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20404 2264 20913 2292
rect 20404 2252 20410 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 24118 2252 24124 2304
rect 24176 2292 24182 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24176 2264 24593 2292
rect 24176 2252 24182 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 26326 2252 26332 2304
rect 26384 2292 26390 2304
rect 27893 2295 27951 2301
rect 27893 2292 27905 2295
rect 26384 2264 27905 2292
rect 26384 2252 26390 2264
rect 27893 2261 27905 2264
rect 27939 2261 27951 2295
rect 27893 2255 27951 2261
rect 30834 2252 30840 2304
rect 30892 2292 30898 2304
rect 33045 2295 33103 2301
rect 33045 2292 33057 2295
rect 30892 2264 33057 2292
rect 30892 2252 30898 2264
rect 33045 2261 33057 2264
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 35621 2295 35679 2301
rect 35621 2292 35633 2295
rect 33192 2264 35633 2292
rect 33192 2252 33198 2264
rect 35621 2261 35633 2264
rect 35667 2261 35679 2295
rect 35621 2255 35679 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 5534 2048 5540 2100
rect 5592 2088 5598 2100
rect 8386 2088 8392 2100
rect 5592 2060 8392 2088
rect 5592 2048 5598 2060
rect 8386 2048 8392 2060
rect 8444 2048 8450 2100
rect 9214 2048 9220 2100
rect 9272 2088 9278 2100
rect 14366 2088 14372 2100
rect 9272 2060 14372 2088
rect 9272 2048 9278 2060
rect 14366 2048 14372 2060
rect 14424 2048 14430 2100
rect 18598 2088 18604 2100
rect 16546 2060 18604 2088
rect 2682 1980 2688 2032
rect 2740 2020 2746 2032
rect 12158 2020 12164 2032
rect 2740 1992 12164 2020
rect 2740 1980 2746 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 2498 1912 2504 1964
rect 2556 1952 2562 1964
rect 2556 1924 2774 1952
rect 2556 1912 2562 1924
rect 2746 1884 2774 1924
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 16546 1952 16574 2060
rect 18598 2048 18604 2060
rect 18656 2048 18662 2100
rect 3844 1924 16574 1952
rect 3844 1912 3850 1924
rect 11422 1884 11428 1896
rect 2746 1856 11428 1884
rect 11422 1844 11428 1856
rect 11480 1844 11486 1896
rect 6086 1776 6092 1828
rect 6144 1816 6150 1828
rect 9490 1816 9496 1828
rect 6144 1788 9496 1816
rect 6144 1776 6150 1788
rect 9490 1776 9496 1788
rect 9548 1776 9554 1828
rect 5166 1708 5172 1760
rect 5224 1748 5230 1760
rect 11238 1748 11244 1760
rect 5224 1720 11244 1748
rect 5224 1708 5230 1720
rect 11238 1708 11244 1720
rect 11296 1708 11302 1760
rect 198 1640 204 1692
rect 256 1680 262 1692
rect 8478 1680 8484 1692
rect 256 1652 8484 1680
rect 256 1640 262 1652
rect 8478 1640 8484 1652
rect 8536 1640 8542 1692
rect 5442 1572 5448 1624
rect 5500 1612 5506 1624
rect 8754 1612 8760 1624
rect 5500 1584 8760 1612
rect 5500 1572 5506 1584
rect 8754 1572 8760 1584
rect 8812 1572 8818 1624
rect 3602 1368 3608 1420
rect 3660 1408 3666 1420
rect 5350 1408 5356 1420
rect 3660 1380 5356 1408
rect 3660 1368 3666 1380
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 6546 1408 6552 1420
rect 6052 1380 6552 1408
rect 6052 1368 6058 1380
rect 6546 1368 6552 1380
rect 6604 1368 6610 1420
rect 6730 1368 6736 1420
rect 6788 1408 6794 1420
rect 9122 1408 9128 1420
rect 6788 1380 9128 1408
rect 6788 1368 6794 1380
rect 9122 1368 9128 1380
rect 9180 1368 9186 1420
rect 1946 1096 1952 1148
rect 2004 1136 2010 1148
rect 6178 1136 6184 1148
rect 2004 1108 6184 1136
rect 2004 1096 2010 1108
rect 6178 1096 6184 1108
rect 6236 1096 6242 1148
rect 10318 1096 10324 1148
rect 10376 1136 10382 1148
rect 11790 1136 11796 1148
rect 10376 1108 11796 1136
rect 10376 1096 10382 1108
rect 11790 1096 11796 1108
rect 11848 1096 11854 1148
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 23572 16600 23624 16652
rect 23020 16532 23072 16584
rect 23756 16532 23808 16584
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 27804 16532 27856 16584
rect 28816 16532 28868 16584
rect 23572 16464 23624 16516
rect 26976 16464 27028 16516
rect 28908 16464 28960 16516
rect 22652 16396 22704 16448
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 26240 16396 26292 16448
rect 27160 16396 27212 16448
rect 28356 16439 28408 16448
rect 28356 16405 28371 16439
rect 28371 16405 28405 16439
rect 28405 16405 28408 16439
rect 28356 16396 28408 16405
rect 29092 16396 29144 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 23572 16192 23624 16244
rect 20720 15988 20772 16040
rect 22652 16099 22704 16108
rect 22652 16065 22686 16099
rect 22686 16065 22704 16099
rect 22652 16056 22704 16065
rect 25136 16124 25188 16176
rect 24308 16056 24360 16108
rect 26240 16056 26292 16108
rect 23480 15920 23532 15972
rect 23848 15852 23900 15904
rect 26700 15988 26752 16040
rect 28356 16056 28408 16108
rect 30288 16056 30340 16108
rect 30748 16056 30800 16108
rect 32496 16056 32548 16108
rect 26976 15963 27028 15972
rect 26976 15929 26985 15963
rect 26985 15929 27019 15963
rect 27019 15929 27028 15963
rect 26976 15920 27028 15929
rect 29000 15852 29052 15904
rect 29184 15852 29236 15904
rect 31300 15852 31352 15904
rect 31576 15895 31628 15904
rect 31576 15861 31585 15895
rect 31585 15861 31619 15895
rect 31619 15861 31628 15895
rect 31576 15852 31628 15861
rect 32128 15895 32180 15904
rect 32128 15861 32137 15895
rect 32137 15861 32171 15895
rect 32171 15861 32180 15895
rect 32128 15852 32180 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 22652 15648 22704 15700
rect 23020 15691 23072 15700
rect 23020 15657 23029 15691
rect 23029 15657 23063 15691
rect 23063 15657 23072 15691
rect 23020 15648 23072 15657
rect 24308 15648 24360 15700
rect 28908 15691 28960 15700
rect 28908 15657 28917 15691
rect 28917 15657 28951 15691
rect 28951 15657 28960 15691
rect 28908 15648 28960 15657
rect 30288 15648 30340 15700
rect 30748 15691 30800 15700
rect 30748 15657 30757 15691
rect 30757 15657 30791 15691
rect 30791 15657 30800 15691
rect 30748 15648 30800 15657
rect 28816 15623 28868 15632
rect 28816 15589 28825 15623
rect 28825 15589 28859 15623
rect 28859 15589 28868 15623
rect 28816 15580 28868 15589
rect 31944 15648 31996 15700
rect 29000 15555 29052 15564
rect 29000 15521 29009 15555
rect 29009 15521 29043 15555
rect 29043 15521 29052 15555
rect 29000 15512 29052 15521
rect 20720 15444 20772 15496
rect 21824 15376 21876 15428
rect 23664 15444 23716 15496
rect 23756 15487 23808 15496
rect 23756 15453 23765 15487
rect 23765 15453 23799 15487
rect 23799 15453 23808 15487
rect 23756 15444 23808 15453
rect 24952 15444 25004 15496
rect 25136 15444 25188 15496
rect 27160 15487 27212 15496
rect 27160 15453 27194 15487
rect 27194 15453 27212 15487
rect 27160 15444 27212 15453
rect 29092 15444 29144 15496
rect 31116 15512 31168 15564
rect 23388 15376 23440 15428
rect 21916 15308 21968 15360
rect 22836 15351 22888 15360
rect 22836 15317 22845 15351
rect 22845 15317 22879 15351
rect 22879 15317 22888 15351
rect 22836 15308 22888 15317
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 30472 15376 30524 15428
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 31300 15487 31352 15496
rect 30656 15444 30708 15453
rect 31300 15453 31309 15487
rect 31309 15453 31343 15487
rect 31343 15453 31352 15487
rect 31300 15444 31352 15453
rect 32128 15444 32180 15496
rect 25596 15308 25648 15360
rect 27896 15308 27948 15360
rect 32312 15308 32364 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 22836 15104 22888 15156
rect 20444 14968 20496 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23020 15036 23072 15088
rect 24952 15104 25004 15156
rect 27804 15147 27856 15156
rect 27804 15113 27813 15147
rect 27813 15113 27847 15147
rect 27847 15113 27856 15147
rect 27804 15104 27856 15113
rect 30656 15104 30708 15156
rect 25412 15079 25464 15088
rect 25412 15045 25421 15079
rect 25421 15045 25455 15079
rect 25455 15045 25464 15079
rect 25412 15036 25464 15045
rect 27344 15036 27396 15088
rect 23848 15011 23900 15020
rect 21916 14900 21968 14952
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 26424 14968 26476 15020
rect 27896 14968 27948 15020
rect 31576 15036 31628 15088
rect 31392 14968 31444 15020
rect 26700 14900 26752 14952
rect 27804 14900 27856 14952
rect 28816 14900 28868 14952
rect 20720 14764 20772 14816
rect 21364 14764 21416 14816
rect 22192 14807 22244 14816
rect 22192 14773 22201 14807
rect 22201 14773 22235 14807
rect 22235 14773 22244 14807
rect 22192 14764 22244 14773
rect 24400 14764 24452 14816
rect 24768 14764 24820 14816
rect 26148 14832 26200 14884
rect 26056 14807 26108 14816
rect 26056 14773 26065 14807
rect 26065 14773 26099 14807
rect 26099 14773 26108 14807
rect 26056 14764 26108 14773
rect 28632 14807 28684 14816
rect 28632 14773 28641 14807
rect 28641 14773 28675 14807
rect 28675 14773 28684 14807
rect 28632 14764 28684 14773
rect 32312 14807 32364 14816
rect 32312 14773 32321 14807
rect 32321 14773 32355 14807
rect 32355 14773 32364 14807
rect 32312 14764 32364 14773
rect 32496 14807 32548 14816
rect 32496 14773 32505 14807
rect 32505 14773 32539 14807
rect 32539 14773 32548 14807
rect 32496 14764 32548 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 17592 14288 17644 14340
rect 20076 14424 20128 14476
rect 20444 14560 20496 14612
rect 22008 14560 22060 14612
rect 23388 14603 23440 14612
rect 23388 14569 23397 14603
rect 23397 14569 23431 14603
rect 23431 14569 23440 14603
rect 23388 14560 23440 14569
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 25412 14603 25464 14612
rect 25412 14569 25421 14603
rect 25421 14569 25455 14603
rect 25455 14569 25464 14603
rect 25412 14560 25464 14569
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 27344 14603 27396 14612
rect 27344 14569 27353 14603
rect 27353 14569 27387 14603
rect 27387 14569 27396 14603
rect 27344 14560 27396 14569
rect 28724 14560 28776 14612
rect 30472 14560 30524 14612
rect 23296 14492 23348 14544
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 21364 14356 21416 14408
rect 25872 14492 25924 14544
rect 31116 14424 31168 14476
rect 22192 14399 22244 14408
rect 22192 14365 22201 14399
rect 22201 14365 22235 14399
rect 22235 14365 22244 14399
rect 23020 14399 23072 14408
rect 22192 14356 22244 14365
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 24308 14356 24360 14408
rect 25044 14356 25096 14408
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 26516 14399 26568 14408
rect 26516 14365 26525 14399
rect 26525 14365 26559 14399
rect 26559 14365 26568 14399
rect 26516 14356 26568 14365
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20260 14263 20312 14272
rect 20260 14229 20269 14263
rect 20269 14229 20303 14263
rect 20303 14229 20312 14263
rect 20260 14220 20312 14229
rect 25136 14288 25188 14340
rect 27712 14356 27764 14408
rect 28632 14356 28684 14408
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 30196 14399 30248 14408
rect 30196 14365 30205 14399
rect 30205 14365 30239 14399
rect 30239 14365 30248 14399
rect 30196 14356 30248 14365
rect 30380 14399 30432 14408
rect 30380 14365 30389 14399
rect 30389 14365 30423 14399
rect 30423 14365 30432 14399
rect 30380 14356 30432 14365
rect 27896 14288 27948 14340
rect 21824 14220 21876 14272
rect 22008 14220 22060 14272
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 25320 14220 25372 14272
rect 27804 14220 27856 14272
rect 27988 14220 28040 14272
rect 28908 14220 28960 14272
rect 29000 14220 29052 14272
rect 29644 14220 29696 14272
rect 31484 14356 31536 14408
rect 31392 14288 31444 14340
rect 31576 14220 31628 14272
rect 31760 14263 31812 14272
rect 31760 14229 31769 14263
rect 31769 14229 31803 14263
rect 31803 14229 31812 14263
rect 31760 14220 31812 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 18604 14016 18656 14068
rect 19248 13948 19300 14000
rect 20444 14016 20496 14068
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 27988 14016 28040 14068
rect 28908 14016 28960 14068
rect 29736 14016 29788 14068
rect 31484 14059 31536 14068
rect 31484 14025 31493 14059
rect 31493 14025 31527 14059
rect 31527 14025 31536 14059
rect 31484 14016 31536 14025
rect 21364 13948 21416 14000
rect 21548 13948 21600 14000
rect 21916 13948 21968 14000
rect 20076 13880 20128 13932
rect 16948 13812 17000 13864
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 22376 13880 22428 13932
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25596 13948 25648 14000
rect 25964 13948 26016 14000
rect 26240 13991 26292 14000
rect 26240 13957 26249 13991
rect 26249 13957 26283 13991
rect 26283 13957 26292 13991
rect 26240 13948 26292 13957
rect 27620 13991 27672 14000
rect 27620 13957 27629 13991
rect 27629 13957 27663 13991
rect 27663 13957 27672 13991
rect 27620 13948 27672 13957
rect 28356 13948 28408 14000
rect 27712 13880 27764 13932
rect 27988 13880 28040 13932
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 28632 13923 28684 13932
rect 28632 13889 28641 13923
rect 28641 13889 28675 13923
rect 28675 13889 28684 13923
rect 28632 13880 28684 13889
rect 29092 13948 29144 14000
rect 31300 13948 31352 14000
rect 31760 13948 31812 14000
rect 21180 13812 21232 13864
rect 21456 13812 21508 13864
rect 22008 13812 22060 13864
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 23020 13855 23072 13864
rect 23020 13821 23029 13855
rect 23029 13821 23063 13855
rect 23063 13821 23072 13855
rect 23020 13812 23072 13821
rect 23664 13812 23716 13864
rect 24492 13812 24544 13864
rect 24860 13812 24912 13864
rect 26516 13812 26568 13864
rect 29644 13923 29696 13932
rect 29644 13889 29678 13923
rect 29678 13889 29696 13923
rect 29644 13880 29696 13889
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 19432 13744 19484 13796
rect 23480 13744 23532 13796
rect 29276 13812 29328 13864
rect 30380 13812 30432 13864
rect 30932 13812 30984 13864
rect 31116 13744 31168 13796
rect 31668 13880 31720 13932
rect 33692 14016 33744 14068
rect 21088 13719 21140 13728
rect 21088 13685 21097 13719
rect 21097 13685 21131 13719
rect 21131 13685 21140 13719
rect 21088 13676 21140 13685
rect 22008 13719 22060 13728
rect 22008 13685 22017 13719
rect 22017 13685 22051 13719
rect 22051 13685 22060 13719
rect 22008 13676 22060 13685
rect 22284 13676 22336 13728
rect 26148 13676 26200 13728
rect 29552 13676 29604 13728
rect 30748 13719 30800 13728
rect 30748 13685 30757 13719
rect 30757 13685 30791 13719
rect 30791 13685 30800 13719
rect 30748 13676 30800 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 22284 13472 22336 13524
rect 32496 13472 32548 13524
rect 14924 13268 14976 13320
rect 20812 13404 20864 13456
rect 20904 13404 20956 13456
rect 21548 13404 21600 13456
rect 29276 13404 29328 13456
rect 30748 13404 30800 13456
rect 20168 13336 20220 13388
rect 20720 13336 20772 13388
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 24952 13336 25004 13388
rect 20076 13268 20128 13320
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21732 13268 21784 13320
rect 19984 13200 20036 13252
rect 17132 13132 17184 13184
rect 19340 13132 19392 13184
rect 19432 13132 19484 13184
rect 20996 13132 21048 13184
rect 22928 13200 22980 13252
rect 22008 13132 22060 13184
rect 22100 13132 22152 13184
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 26148 13336 26200 13388
rect 29552 13379 29604 13388
rect 29552 13345 29561 13379
rect 29561 13345 29595 13379
rect 29595 13345 29604 13379
rect 29552 13336 29604 13345
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 31944 13336 31996 13388
rect 24860 13268 24912 13277
rect 25044 13200 25096 13252
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 27528 13311 27580 13320
rect 26516 13268 26568 13277
rect 27528 13277 27537 13311
rect 27537 13277 27571 13311
rect 27571 13277 27580 13311
rect 27528 13268 27580 13277
rect 29000 13268 29052 13320
rect 31208 13268 31260 13320
rect 32404 13268 32456 13320
rect 30288 13200 30340 13252
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 26332 13175 26384 13184
rect 26332 13141 26341 13175
rect 26341 13141 26375 13175
rect 26375 13141 26384 13175
rect 26332 13132 26384 13141
rect 26424 13132 26476 13184
rect 27344 13132 27396 13184
rect 28448 13132 28500 13184
rect 28724 13132 28776 13184
rect 31208 13175 31260 13184
rect 31208 13141 31217 13175
rect 31217 13141 31251 13175
rect 31251 13141 31260 13175
rect 31392 13175 31444 13184
rect 31208 13132 31260 13141
rect 31392 13141 31401 13175
rect 31401 13141 31435 13175
rect 31435 13141 31444 13175
rect 31392 13132 31444 13141
rect 31484 13132 31536 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 20996 12928 21048 12980
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 22376 12928 22428 12937
rect 24216 12928 24268 12980
rect 24584 12928 24636 12980
rect 19248 12903 19300 12912
rect 19248 12869 19257 12903
rect 19257 12869 19291 12903
rect 19291 12869 19300 12903
rect 19248 12860 19300 12869
rect 26240 12928 26292 12980
rect 27620 12928 27672 12980
rect 30932 12971 30984 12980
rect 9680 12835 9732 12844
rect 9680 12801 9697 12835
rect 9697 12801 9731 12835
rect 9731 12801 9732 12835
rect 10508 12835 10560 12844
rect 9680 12792 9732 12801
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 17684 12792 17736 12844
rect 19432 12792 19484 12844
rect 19984 12792 20036 12844
rect 21640 12792 21692 12844
rect 25320 12835 25372 12844
rect 25320 12801 25329 12835
rect 25329 12801 25363 12835
rect 25363 12801 25372 12835
rect 25320 12792 25372 12801
rect 20260 12724 20312 12776
rect 22284 12724 22336 12776
rect 17592 12656 17644 12708
rect 17960 12656 18012 12708
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 11612 12588 11664 12640
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 19156 12588 19208 12640
rect 20812 12588 20864 12640
rect 22652 12588 22704 12640
rect 26148 12835 26200 12844
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 26424 12792 26476 12844
rect 26976 12792 27028 12844
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 28632 12792 28684 12844
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 26332 12767 26384 12776
rect 26332 12733 26341 12767
rect 26341 12733 26375 12767
rect 26375 12733 26384 12767
rect 26332 12724 26384 12733
rect 26884 12724 26936 12776
rect 27988 12724 28040 12776
rect 28356 12724 28408 12776
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 30656 12860 30708 12912
rect 30932 12937 30941 12971
rect 30941 12937 30975 12971
rect 30975 12937 30984 12971
rect 30932 12928 30984 12937
rect 31392 12928 31444 12980
rect 31024 12860 31076 12912
rect 31208 12860 31260 12912
rect 31300 12792 31352 12844
rect 31484 12792 31536 12844
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 32404 12835 32456 12844
rect 32404 12801 32413 12835
rect 32413 12801 32447 12835
rect 32447 12801 32456 12835
rect 32404 12792 32456 12801
rect 33140 12792 33192 12844
rect 26516 12656 26568 12708
rect 28080 12656 28132 12708
rect 28724 12656 28776 12708
rect 29000 12588 29052 12640
rect 29644 12588 29696 12640
rect 29920 12588 29972 12640
rect 30288 12588 30340 12640
rect 31392 12631 31444 12640
rect 31392 12597 31401 12631
rect 31401 12597 31435 12631
rect 31435 12597 31444 12631
rect 31392 12588 31444 12597
rect 33324 12724 33376 12776
rect 33876 12767 33928 12776
rect 31576 12656 31628 12708
rect 33508 12656 33560 12708
rect 33876 12733 33885 12767
rect 33885 12733 33919 12767
rect 33919 12733 33928 12767
rect 33876 12724 33928 12733
rect 32220 12588 32272 12640
rect 32680 12631 32732 12640
rect 32680 12597 32689 12631
rect 32689 12597 32723 12631
rect 32723 12597 32732 12631
rect 32680 12588 32732 12597
rect 33968 12588 34020 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10508 12384 10560 12436
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 19156 12384 19208 12436
rect 19984 12384 20036 12436
rect 18420 12316 18472 12368
rect 8300 12248 8352 12300
rect 9496 12248 9548 12300
rect 18052 12248 18104 12300
rect 21732 12384 21784 12436
rect 24768 12384 24820 12436
rect 24952 12384 25004 12436
rect 24492 12316 24544 12368
rect 23296 12291 23348 12300
rect 23296 12257 23305 12291
rect 23305 12257 23339 12291
rect 23339 12257 23348 12291
rect 23296 12248 23348 12257
rect 24400 12248 24452 12300
rect 27160 12316 27212 12368
rect 30196 12384 30248 12436
rect 31116 12248 31168 12300
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 8576 12180 8628 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 13820 12180 13872 12232
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 9956 12112 10008 12164
rect 10508 12155 10560 12164
rect 10508 12121 10517 12155
rect 10517 12121 10551 12155
rect 10551 12121 10560 12155
rect 10508 12112 10560 12121
rect 14832 12112 14884 12164
rect 5816 12044 5868 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 9220 12044 9272 12096
rect 10416 12044 10468 12096
rect 10692 12044 10744 12096
rect 12440 12044 12492 12096
rect 19156 12180 19208 12232
rect 20720 12180 20772 12232
rect 21364 12180 21416 12232
rect 21640 12180 21692 12232
rect 21732 12180 21784 12232
rect 17500 12112 17552 12164
rect 20076 12112 20128 12164
rect 20536 12112 20588 12164
rect 21088 12112 21140 12164
rect 21180 12112 21232 12164
rect 17408 12044 17460 12096
rect 19432 12044 19484 12096
rect 21364 12044 21416 12096
rect 21548 12044 21600 12096
rect 21824 12044 21876 12096
rect 22376 12112 22428 12164
rect 22744 12112 22796 12164
rect 25596 12223 25648 12232
rect 24584 12112 24636 12164
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 27712 12223 27764 12232
rect 27712 12189 27721 12223
rect 27721 12189 27755 12223
rect 27755 12189 27764 12223
rect 27712 12180 27764 12189
rect 27988 12180 28040 12232
rect 26056 12112 26108 12164
rect 25688 12044 25740 12096
rect 28632 12155 28684 12164
rect 26976 12087 27028 12096
rect 26976 12053 26985 12087
rect 26985 12053 27019 12087
rect 27019 12053 27028 12087
rect 26976 12044 27028 12053
rect 27804 12044 27856 12096
rect 28264 12044 28316 12096
rect 28632 12121 28641 12155
rect 28641 12121 28675 12155
rect 28675 12121 28684 12155
rect 28632 12112 28684 12121
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 30748 12223 30800 12232
rect 29920 12180 29972 12189
rect 30748 12189 30757 12223
rect 30757 12189 30791 12223
rect 30791 12189 30800 12223
rect 30748 12180 30800 12189
rect 31208 12223 31260 12232
rect 31208 12189 31217 12223
rect 31217 12189 31251 12223
rect 31251 12189 31260 12223
rect 31208 12180 31260 12189
rect 32680 12180 32732 12232
rect 33324 12223 33376 12232
rect 33324 12189 33333 12223
rect 33333 12189 33367 12223
rect 33367 12189 33376 12223
rect 33324 12180 33376 12189
rect 30656 12112 30708 12164
rect 31484 12155 31536 12164
rect 31484 12121 31518 12155
rect 31518 12121 31536 12155
rect 31484 12112 31536 12121
rect 31668 12112 31720 12164
rect 29644 12044 29696 12096
rect 30564 12087 30616 12096
rect 30564 12053 30573 12087
rect 30573 12053 30607 12087
rect 30607 12053 30616 12087
rect 30564 12044 30616 12053
rect 32588 12087 32640 12096
rect 32588 12053 32597 12087
rect 32597 12053 32631 12087
rect 32631 12053 32640 12087
rect 32588 12044 32640 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 12532 11840 12584 11892
rect 21180 11840 21232 11892
rect 22008 11840 22060 11892
rect 22376 11883 22428 11892
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 22928 11883 22980 11892
rect 22928 11849 22937 11883
rect 22937 11849 22971 11883
rect 22971 11849 22980 11883
rect 22928 11840 22980 11849
rect 29000 11840 29052 11892
rect 31024 11883 31076 11892
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 7012 11772 7064 11824
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 10416 11772 10468 11824
rect 11612 11772 11664 11824
rect 13268 11772 13320 11824
rect 9220 11704 9272 11756
rect 12348 11704 12400 11756
rect 13360 11747 13412 11756
rect 13360 11713 13369 11747
rect 13369 11713 13403 11747
rect 13403 11713 13412 11747
rect 13360 11704 13412 11713
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14556 11704 14608 11756
rect 15108 11704 15160 11756
rect 8300 11636 8352 11688
rect 17500 11704 17552 11756
rect 20720 11772 20772 11824
rect 22284 11772 22336 11824
rect 20536 11704 20588 11756
rect 22100 11704 22152 11756
rect 23020 11747 23072 11756
rect 16672 11636 16724 11688
rect 16764 11636 16816 11688
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 21916 11636 21968 11688
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 25596 11772 25648 11824
rect 26608 11772 26660 11824
rect 24676 11747 24728 11756
rect 24676 11713 24710 11747
rect 24710 11713 24728 11747
rect 26424 11747 26476 11756
rect 24676 11704 24728 11713
rect 26424 11713 26433 11747
rect 26433 11713 26467 11747
rect 26467 11713 26476 11747
rect 26424 11704 26476 11713
rect 27528 11772 27580 11824
rect 30564 11772 30616 11824
rect 27068 11704 27120 11756
rect 31024 11849 31033 11883
rect 31033 11849 31067 11883
rect 31067 11849 31076 11883
rect 31024 11840 31076 11849
rect 31668 11772 31720 11824
rect 23756 11636 23808 11688
rect 16856 11568 16908 11620
rect 18604 11568 18656 11620
rect 21824 11611 21876 11620
rect 6736 11500 6788 11552
rect 10324 11500 10376 11552
rect 13268 11500 13320 11552
rect 14188 11500 14240 11552
rect 14464 11500 14516 11552
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 18144 11500 18196 11552
rect 19156 11500 19208 11552
rect 21364 11500 21416 11552
rect 21824 11577 21833 11611
rect 21833 11577 21867 11611
rect 21867 11577 21876 11611
rect 21824 11568 21876 11577
rect 22008 11568 22060 11620
rect 22560 11500 22612 11552
rect 26884 11568 26936 11620
rect 25780 11543 25832 11552
rect 25780 11509 25789 11543
rect 25789 11509 25823 11543
rect 25823 11509 25832 11543
rect 26240 11543 26292 11552
rect 25780 11500 25832 11509
rect 26240 11509 26249 11543
rect 26249 11509 26283 11543
rect 26283 11509 26292 11543
rect 26240 11500 26292 11509
rect 28264 11500 28316 11552
rect 32772 11704 32824 11756
rect 30932 11636 30984 11688
rect 32956 11636 33008 11688
rect 29552 11500 29604 11552
rect 31208 11568 31260 11620
rect 34152 11636 34204 11688
rect 33324 11500 33376 11552
rect 34428 11543 34480 11552
rect 34428 11509 34437 11543
rect 34437 11509 34471 11543
rect 34471 11509 34480 11543
rect 34428 11500 34480 11509
rect 36268 11543 36320 11552
rect 36268 11509 36277 11543
rect 36277 11509 36311 11543
rect 36311 11509 36320 11543
rect 36268 11500 36320 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7748 11296 7800 11348
rect 12532 11296 12584 11348
rect 12716 11296 12768 11348
rect 14004 11296 14056 11348
rect 15752 11296 15804 11348
rect 16672 11296 16724 11348
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 23664 11296 23716 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 25044 11339 25096 11348
rect 25044 11305 25053 11339
rect 25053 11305 25087 11339
rect 25087 11305 25096 11339
rect 25044 11296 25096 11305
rect 25872 11296 25924 11348
rect 27068 11296 27120 11348
rect 27712 11296 27764 11348
rect 28632 11296 28684 11348
rect 30748 11296 30800 11348
rect 34152 11296 34204 11348
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 9680 11160 9732 11212
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 7656 11092 7708 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 14832 11228 14884 11280
rect 18236 11228 18288 11280
rect 24308 11228 24360 11280
rect 26884 11228 26936 11280
rect 33876 11228 33928 11280
rect 12624 11160 12676 11212
rect 13268 11160 13320 11212
rect 18144 11160 18196 11212
rect 18420 11203 18472 11212
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 5632 11024 5684 11076
rect 10692 11067 10744 11076
rect 10692 11033 10726 11067
rect 10726 11033 10744 11067
rect 10692 11024 10744 11033
rect 13176 11024 13228 11076
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 11428 10956 11480 11008
rect 12348 10956 12400 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 15292 11024 15344 11076
rect 18052 11092 18104 11144
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 19984 11160 20036 11212
rect 16764 11024 16816 11076
rect 17960 11024 18012 11076
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 18604 11092 18656 11144
rect 19432 11092 19484 11144
rect 20812 11092 20864 11144
rect 22376 11160 22428 11212
rect 22192 11092 22244 11144
rect 20904 11024 20956 11076
rect 23020 11092 23072 11144
rect 26148 11160 26200 11212
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 23204 11024 23256 11076
rect 16488 10999 16540 11008
rect 16488 10965 16497 10999
rect 16497 10965 16531 10999
rect 16531 10965 16540 10999
rect 16488 10956 16540 10965
rect 17684 10956 17736 11008
rect 25320 11024 25372 11076
rect 25044 10956 25096 11008
rect 25688 11024 25740 11076
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 28264 11160 28316 11212
rect 29920 11160 29972 11212
rect 27160 11135 27212 11144
rect 27160 11101 27169 11135
rect 27169 11101 27203 11135
rect 27203 11101 27212 11135
rect 27160 11092 27212 11101
rect 27344 11092 27396 11144
rect 28908 11092 28960 11144
rect 29828 11092 29880 11144
rect 32680 11203 32732 11212
rect 32680 11169 32689 11203
rect 32689 11169 32723 11203
rect 32723 11169 32732 11203
rect 32680 11160 32732 11169
rect 30656 11092 30708 11144
rect 31024 11135 31076 11144
rect 25780 10999 25832 11008
rect 25780 10965 25789 10999
rect 25789 10965 25823 10999
rect 25823 10965 25832 10999
rect 25780 10956 25832 10965
rect 25872 10956 25924 11008
rect 27344 10956 27396 11008
rect 31024 11101 31033 11135
rect 31033 11101 31067 11135
rect 31067 11101 31076 11135
rect 31024 11092 31076 11101
rect 33508 11092 33560 11144
rect 33968 11135 34020 11144
rect 33968 11101 33977 11135
rect 33977 11101 34011 11135
rect 34011 11101 34020 11135
rect 33968 11092 34020 11101
rect 34152 11135 34204 11144
rect 34152 11101 34161 11135
rect 34161 11101 34195 11135
rect 34195 11101 34204 11135
rect 34152 11092 34204 11101
rect 30564 10999 30616 11008
rect 30564 10965 30573 10999
rect 30573 10965 30607 10999
rect 30607 10965 30616 10999
rect 30564 10956 30616 10965
rect 30932 10956 30984 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 6920 10752 6972 10804
rect 8300 10752 8352 10804
rect 9588 10752 9640 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 11336 10752 11388 10804
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 2412 10548 2464 10600
rect 7196 10616 7248 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 10324 10684 10376 10736
rect 12440 10684 12492 10736
rect 12716 10684 12768 10736
rect 17684 10795 17736 10804
rect 14004 10684 14056 10736
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 8300 10548 8352 10600
rect 3240 10480 3292 10532
rect 9312 10616 9364 10668
rect 10600 10659 10652 10668
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11428 10616 11480 10668
rect 12348 10659 12400 10668
rect 12348 10625 12357 10659
rect 12357 10625 12391 10659
rect 12391 10625 12400 10659
rect 12348 10616 12400 10625
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 18512 10752 18564 10804
rect 19248 10752 19300 10804
rect 14832 10684 14884 10736
rect 17408 10684 17460 10736
rect 18144 10684 18196 10736
rect 18420 10684 18472 10736
rect 14372 10616 14424 10668
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 14280 10548 14332 10600
rect 15108 10548 15160 10600
rect 15844 10548 15896 10600
rect 16948 10616 17000 10668
rect 18052 10616 18104 10668
rect 21364 10684 21416 10736
rect 21456 10684 21508 10736
rect 22836 10752 22888 10804
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 23572 10684 23624 10736
rect 22100 10616 22152 10668
rect 23112 10616 23164 10668
rect 23940 10684 23992 10736
rect 23848 10659 23900 10668
rect 23848 10625 23857 10659
rect 23857 10625 23891 10659
rect 23891 10625 23900 10659
rect 23848 10616 23900 10625
rect 24676 10616 24728 10668
rect 25596 10659 25648 10668
rect 25596 10625 25605 10659
rect 25605 10625 25639 10659
rect 25639 10625 25648 10659
rect 25596 10616 25648 10625
rect 28356 10752 28408 10804
rect 30932 10795 30984 10804
rect 17500 10523 17552 10532
rect 2872 10412 2924 10464
rect 9496 10412 9548 10464
rect 15384 10412 15436 10464
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 18512 10523 18564 10532
rect 18512 10489 18521 10523
rect 18521 10489 18555 10523
rect 18555 10489 18564 10523
rect 18512 10480 18564 10489
rect 19156 10591 19208 10600
rect 19156 10557 19165 10591
rect 19165 10557 19199 10591
rect 19199 10557 19208 10591
rect 19156 10548 19208 10557
rect 19892 10548 19944 10600
rect 20352 10523 20404 10532
rect 20352 10489 20361 10523
rect 20361 10489 20395 10523
rect 20395 10489 20404 10523
rect 20352 10480 20404 10489
rect 22468 10480 22520 10532
rect 24216 10480 24268 10532
rect 16580 10412 16632 10464
rect 16948 10412 17000 10464
rect 19892 10412 19944 10464
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 22928 10412 22980 10464
rect 23204 10412 23256 10464
rect 23480 10455 23532 10464
rect 23480 10421 23489 10455
rect 23489 10421 23523 10455
rect 23523 10421 23532 10455
rect 23480 10412 23532 10421
rect 25504 10412 25556 10464
rect 25688 10412 25740 10464
rect 28448 10684 28500 10736
rect 30564 10684 30616 10736
rect 30932 10761 30941 10795
rect 30941 10761 30975 10795
rect 30975 10761 30984 10795
rect 30932 10752 30984 10761
rect 33140 10752 33192 10804
rect 34244 10752 34296 10804
rect 31392 10684 31444 10736
rect 26516 10616 26568 10668
rect 28908 10659 28960 10668
rect 28908 10625 28917 10659
rect 28917 10625 28951 10659
rect 28951 10625 28960 10659
rect 28908 10616 28960 10625
rect 29552 10659 29604 10668
rect 29552 10625 29561 10659
rect 29561 10625 29595 10659
rect 29595 10625 29604 10659
rect 29552 10616 29604 10625
rect 29644 10616 29696 10668
rect 30932 10616 30984 10668
rect 31668 10616 31720 10668
rect 33324 10684 33376 10736
rect 33416 10616 33468 10668
rect 34428 10616 34480 10668
rect 33324 10548 33376 10600
rect 29092 10523 29144 10532
rect 26608 10412 26660 10464
rect 29092 10489 29101 10523
rect 29101 10489 29135 10523
rect 29135 10489 29144 10523
rect 29092 10480 29144 10489
rect 30564 10480 30616 10532
rect 32772 10523 32824 10532
rect 30748 10412 30800 10464
rect 30840 10412 30892 10464
rect 31944 10412 31996 10464
rect 32772 10489 32781 10523
rect 32781 10489 32815 10523
rect 32815 10489 32824 10523
rect 32772 10480 32824 10489
rect 34152 10480 34204 10532
rect 34612 10412 34664 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 7932 10208 7984 10260
rect 8392 10208 8444 10260
rect 9772 10208 9824 10260
rect 11060 10208 11112 10260
rect 12164 10208 12216 10260
rect 4712 10140 4764 10192
rect 7196 10140 7248 10192
rect 6184 10004 6236 10056
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 5356 9936 5408 9988
rect 5816 9936 5868 9988
rect 7196 10004 7248 10056
rect 7748 10004 7800 10056
rect 10508 10140 10560 10192
rect 15384 10208 15436 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 17960 10208 18012 10260
rect 18604 10208 18656 10260
rect 21180 10208 21232 10260
rect 18328 10183 18380 10192
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11336 10047 11388 10056
rect 6368 9868 6420 9920
rect 6920 9868 6972 9920
rect 8760 9868 8812 9920
rect 9496 9936 9548 9988
rect 10140 9979 10192 9988
rect 10140 9945 10149 9979
rect 10149 9945 10183 9979
rect 10183 9945 10192 9979
rect 10140 9936 10192 9945
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11980 10004 12032 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 14188 10004 14240 10056
rect 18328 10149 18337 10183
rect 18337 10149 18371 10183
rect 18371 10149 18380 10183
rect 18328 10140 18380 10149
rect 18788 10140 18840 10192
rect 28908 10208 28960 10260
rect 30656 10208 30708 10260
rect 31392 10208 31444 10260
rect 32956 10208 33008 10260
rect 33416 10208 33468 10260
rect 28448 10183 28500 10192
rect 15016 10072 15068 10124
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 14556 10004 14608 10056
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 11520 9868 11572 9920
rect 11612 9868 11664 9920
rect 15108 9936 15160 9988
rect 15844 10004 15896 10056
rect 16396 10004 16448 10056
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 16396 9868 16448 9920
rect 17960 9936 18012 9988
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 23020 10004 23072 10056
rect 24584 10047 24636 10056
rect 24584 10013 24591 10047
rect 24591 10013 24636 10047
rect 18052 9868 18104 9920
rect 18420 9868 18472 9920
rect 22652 9936 22704 9988
rect 23756 9936 23808 9988
rect 24584 10004 24636 10013
rect 25596 10072 25648 10124
rect 28448 10149 28457 10183
rect 28457 10149 28491 10183
rect 28491 10149 28500 10183
rect 28448 10140 28500 10149
rect 31208 10140 31260 10192
rect 26608 10115 26660 10124
rect 24860 10004 24912 10056
rect 25320 10004 25372 10056
rect 26608 10081 26617 10115
rect 26617 10081 26651 10115
rect 26651 10081 26660 10115
rect 26608 10072 26660 10081
rect 25412 9936 25464 9988
rect 24952 9868 25004 9920
rect 25044 9911 25096 9920
rect 25044 9877 25053 9911
rect 25053 9877 25087 9911
rect 25087 9877 25096 9911
rect 25872 10004 25924 10056
rect 30840 10072 30892 10124
rect 32496 10072 32548 10124
rect 32956 10072 33008 10124
rect 33508 10115 33560 10124
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28632 10047 28684 10056
rect 28448 10004 28500 10013
rect 28632 10013 28641 10047
rect 28641 10013 28675 10047
rect 28675 10013 28684 10047
rect 28632 10004 28684 10013
rect 29828 10004 29880 10056
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 25044 9868 25096 9877
rect 26056 9868 26108 9920
rect 28448 9868 28500 9920
rect 29644 9936 29696 9988
rect 32128 10004 32180 10056
rect 32404 10047 32456 10056
rect 32404 10013 32413 10047
rect 32413 10013 32447 10047
rect 32447 10013 32456 10047
rect 32404 10004 32456 10013
rect 33048 10047 33100 10056
rect 33048 10013 33057 10047
rect 33057 10013 33091 10047
rect 33091 10013 33100 10047
rect 33048 10004 33100 10013
rect 33232 10004 33284 10056
rect 33508 10081 33517 10115
rect 33517 10081 33551 10115
rect 33551 10081 33560 10115
rect 33508 10072 33560 10081
rect 34152 10047 34204 10056
rect 34152 10013 34161 10047
rect 34161 10013 34195 10047
rect 34195 10013 34204 10047
rect 34152 10004 34204 10013
rect 34428 10004 34480 10056
rect 32036 9936 32088 9988
rect 30656 9868 30708 9920
rect 31024 9868 31076 9920
rect 32220 9911 32272 9920
rect 32220 9877 32229 9911
rect 32229 9877 32263 9911
rect 32263 9877 32272 9911
rect 32220 9868 32272 9877
rect 33140 9868 33192 9920
rect 33784 9936 33836 9988
rect 36268 10004 36320 10056
rect 33600 9868 33652 9920
rect 34060 9911 34112 9920
rect 34060 9877 34069 9911
rect 34069 9877 34103 9911
rect 34103 9877 34112 9911
rect 34060 9868 34112 9877
rect 35624 9868 35676 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2228 9664 2280 9716
rect 11336 9664 11388 9716
rect 11612 9664 11664 9716
rect 16396 9664 16448 9716
rect 16672 9664 16724 9716
rect 20720 9664 20772 9716
rect 21824 9664 21876 9716
rect 23756 9664 23808 9716
rect 24676 9664 24728 9716
rect 25412 9707 25464 9716
rect 25412 9673 25421 9707
rect 25421 9673 25455 9707
rect 25455 9673 25464 9707
rect 25412 9664 25464 9673
rect 25596 9664 25648 9716
rect 2136 9596 2188 9648
rect 4068 9596 4120 9648
rect 4896 9596 4948 9648
rect 7012 9596 7064 9648
rect 5632 9528 5684 9580
rect 5724 9528 5776 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6736 9528 6788 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 9312 9528 9364 9580
rect 10416 9528 10468 9580
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 16580 9596 16632 9648
rect 8392 9460 8444 9512
rect 9680 9460 9732 9512
rect 11796 9460 11848 9512
rect 13544 9528 13596 9580
rect 14464 9528 14516 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 15292 9460 15344 9512
rect 15844 9460 15896 9512
rect 16488 9528 16540 9580
rect 18052 9596 18104 9648
rect 18236 9639 18288 9648
rect 18236 9605 18270 9639
rect 18270 9605 18288 9639
rect 18236 9596 18288 9605
rect 22100 9596 22152 9648
rect 22744 9596 22796 9648
rect 24308 9639 24360 9648
rect 24308 9605 24342 9639
rect 24342 9605 24360 9639
rect 24308 9596 24360 9605
rect 29460 9664 29512 9716
rect 31668 9664 31720 9716
rect 33508 9664 33560 9716
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 17316 9528 17368 9580
rect 17224 9460 17276 9512
rect 17868 9460 17920 9512
rect 20444 9528 20496 9580
rect 20720 9528 20772 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 22284 9528 22336 9580
rect 22468 9571 22520 9580
rect 22468 9537 22502 9571
rect 22502 9537 22520 9571
rect 24032 9571 24084 9580
rect 22468 9528 22520 9537
rect 24032 9537 24041 9571
rect 24041 9537 24075 9571
rect 24075 9537 24084 9571
rect 24032 9528 24084 9537
rect 26792 9596 26844 9648
rect 29092 9596 29144 9648
rect 23756 9460 23808 9512
rect 24860 9528 24912 9580
rect 25872 9571 25924 9580
rect 25872 9537 25881 9571
rect 25881 9537 25915 9571
rect 25915 9537 25924 9571
rect 25872 9528 25924 9537
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 25228 9460 25280 9512
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 31024 9528 31076 9580
rect 31576 9571 31628 9580
rect 26608 9460 26660 9512
rect 6460 9324 6512 9376
rect 7932 9324 7984 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 11980 9324 12032 9376
rect 12164 9324 12216 9376
rect 15384 9324 15436 9376
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 19708 9392 19760 9444
rect 19984 9392 20036 9444
rect 20628 9392 20680 9444
rect 21088 9435 21140 9444
rect 21088 9401 21097 9435
rect 21097 9401 21131 9435
rect 21131 9401 21140 9435
rect 21088 9392 21140 9401
rect 28724 9392 28776 9444
rect 31576 9537 31585 9571
rect 31585 9537 31619 9571
rect 31619 9537 31628 9571
rect 31576 9528 31628 9537
rect 32220 9596 32272 9648
rect 34612 9596 34664 9648
rect 34244 9571 34296 9580
rect 34244 9537 34253 9571
rect 34253 9537 34287 9571
rect 34287 9537 34296 9571
rect 34244 9528 34296 9537
rect 31852 9460 31904 9512
rect 33876 9460 33928 9512
rect 35624 9528 35676 9580
rect 35992 9571 36044 9580
rect 34612 9503 34664 9512
rect 34612 9469 34621 9503
rect 34621 9469 34655 9503
rect 34655 9469 34664 9503
rect 34612 9460 34664 9469
rect 35440 9460 35492 9512
rect 35992 9537 36001 9571
rect 36001 9537 36035 9571
rect 36035 9537 36044 9571
rect 35992 9528 36044 9537
rect 34796 9392 34848 9444
rect 19432 9324 19484 9376
rect 21916 9324 21968 9376
rect 25412 9324 25464 9376
rect 29184 9324 29236 9376
rect 29644 9324 29696 9376
rect 31116 9324 31168 9376
rect 31760 9324 31812 9376
rect 33048 9324 33100 9376
rect 33876 9324 33928 9376
rect 34152 9324 34204 9376
rect 34520 9324 34572 9376
rect 35808 9367 35860 9376
rect 35808 9333 35817 9367
rect 35817 9333 35851 9367
rect 35851 9333 35860 9367
rect 35808 9324 35860 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4068 9120 4120 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 10416 9120 10468 9172
rect 10600 9163 10652 9172
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 12072 9120 12124 9172
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 9036 9052 9088 9104
rect 15292 9120 15344 9172
rect 15384 9120 15436 9172
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 4896 8916 4948 8968
rect 6276 8916 6328 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 4620 8891 4672 8900
rect 4620 8857 4654 8891
rect 4654 8857 4672 8891
rect 4620 8848 4672 8857
rect 5448 8848 5500 8900
rect 7472 8916 7524 8968
rect 7748 8984 7800 9036
rect 8760 8984 8812 9036
rect 11060 9027 11112 9036
rect 6828 8848 6880 8900
rect 8576 8916 8628 8968
rect 8944 8916 8996 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11060 8984 11112 8993
rect 11336 8984 11388 9036
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 9772 8780 9824 8832
rect 11244 8916 11296 8968
rect 11520 8916 11572 8968
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 11428 8848 11480 8900
rect 11980 8916 12032 8968
rect 10968 8780 11020 8832
rect 12072 8780 12124 8832
rect 12348 8780 12400 8832
rect 12532 8780 12584 8832
rect 12900 8848 12952 8900
rect 15752 9052 15804 9104
rect 18880 9120 18932 9172
rect 20168 9120 20220 9172
rect 20812 9120 20864 9172
rect 18328 9052 18380 9104
rect 13360 8984 13412 9036
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 15844 8916 15896 8968
rect 16764 8916 16816 8968
rect 17868 8916 17920 8968
rect 19156 8916 19208 8968
rect 19616 8984 19668 9036
rect 20996 9052 21048 9104
rect 23572 9120 23624 9172
rect 24768 9120 24820 9172
rect 26332 9120 26384 9172
rect 28816 9120 28868 9172
rect 31760 9120 31812 9172
rect 32036 9163 32088 9172
rect 32036 9129 32045 9163
rect 32045 9129 32079 9163
rect 32079 9129 32088 9163
rect 32036 9120 32088 9129
rect 32404 9120 32456 9172
rect 33600 9120 33652 9172
rect 34612 9120 34664 9172
rect 24860 9052 24912 9104
rect 28172 9052 28224 9104
rect 28724 9095 28776 9104
rect 28724 9061 28733 9095
rect 28733 9061 28767 9095
rect 28767 9061 28776 9095
rect 28724 9052 28776 9061
rect 33048 9052 33100 9104
rect 33324 9052 33376 9104
rect 33416 9052 33468 9104
rect 35808 9120 35860 9172
rect 19984 8916 20036 8968
rect 20168 8916 20220 8968
rect 21088 8984 21140 9036
rect 22284 9027 22336 9036
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 21272 8916 21324 8968
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 15752 8780 15804 8832
rect 17592 8780 17644 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19892 8848 19944 8900
rect 20444 8848 20496 8900
rect 22284 8993 22293 9027
rect 22293 8993 22327 9027
rect 22327 8993 22336 9027
rect 22284 8984 22336 8993
rect 24032 8984 24084 9036
rect 26148 8984 26200 9036
rect 26792 9027 26844 9036
rect 26792 8993 26801 9027
rect 26801 8993 26835 9027
rect 26835 8993 26844 9027
rect 26792 8984 26844 8993
rect 29644 9027 29696 9036
rect 26700 8916 26752 8968
rect 22284 8848 22336 8900
rect 22560 8891 22612 8900
rect 22560 8857 22594 8891
rect 22594 8857 22612 8891
rect 22560 8848 22612 8857
rect 22744 8848 22796 8900
rect 27528 8916 27580 8968
rect 28264 8959 28316 8968
rect 28264 8925 28271 8959
rect 28271 8925 28316 8959
rect 28264 8916 28316 8925
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 29644 8993 29653 9027
rect 29653 8993 29687 9027
rect 29687 8993 29696 9027
rect 29644 8984 29696 8993
rect 34060 8984 34112 9036
rect 32220 8916 32272 8968
rect 33232 8916 33284 8968
rect 33508 8916 33560 8968
rect 19432 8780 19484 8832
rect 20352 8780 20404 8832
rect 22376 8780 22428 8832
rect 25228 8780 25280 8832
rect 25320 8780 25372 8832
rect 25872 8780 25924 8832
rect 25964 8780 26016 8832
rect 28908 8848 28960 8900
rect 30748 8848 30800 8900
rect 32312 8848 32364 8900
rect 34520 8916 34572 8968
rect 34704 8959 34756 8968
rect 34704 8925 34713 8959
rect 34713 8925 34747 8959
rect 34747 8925 34756 8959
rect 34704 8916 34756 8925
rect 30472 8780 30524 8832
rect 33784 8891 33836 8900
rect 33784 8857 33793 8891
rect 33793 8857 33827 8891
rect 33827 8857 33836 8891
rect 33784 8848 33836 8857
rect 33968 8891 34020 8900
rect 33968 8857 33993 8891
rect 33993 8857 34020 8891
rect 33968 8848 34020 8857
rect 34428 8848 34480 8900
rect 32680 8823 32732 8832
rect 32680 8789 32689 8823
rect 32689 8789 32723 8823
rect 32723 8789 32732 8823
rect 32680 8780 32732 8789
rect 33140 8823 33192 8832
rect 33140 8789 33149 8823
rect 33149 8789 33183 8823
rect 33183 8789 33192 8823
rect 33140 8780 33192 8789
rect 33600 8780 33652 8832
rect 34796 8780 34848 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 5632 8576 5684 8628
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 9220 8576 9272 8628
rect 16304 8576 16356 8628
rect 16948 8576 17000 8628
rect 20168 8576 20220 8628
rect 21732 8576 21784 8628
rect 6276 8508 6328 8560
rect 6736 8508 6788 8560
rect 9772 8508 9824 8560
rect 10508 8508 10560 8560
rect 5724 8440 5776 8492
rect 5080 8372 5132 8424
rect 6368 8440 6420 8492
rect 7012 8440 7064 8492
rect 7840 8483 7892 8492
rect 7840 8449 7874 8483
rect 7874 8449 7892 8483
rect 9404 8483 9456 8492
rect 7840 8440 7892 8449
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 5540 8304 5592 8356
rect 6644 8304 6696 8356
rect 11336 8372 11388 8424
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 5356 8236 5408 8288
rect 7288 8236 7340 8288
rect 8668 8304 8720 8356
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 13728 8508 13780 8560
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 13544 8372 13596 8424
rect 15476 8440 15528 8492
rect 16488 8440 16540 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17960 8440 18012 8492
rect 19340 8508 19392 8560
rect 19892 8508 19944 8560
rect 22468 8508 22520 8560
rect 22836 8508 22888 8560
rect 19984 8440 20036 8492
rect 20444 8440 20496 8492
rect 16672 8372 16724 8424
rect 13820 8304 13872 8356
rect 14832 8347 14884 8356
rect 14832 8313 14841 8347
rect 14841 8313 14875 8347
rect 14875 8313 14884 8347
rect 14832 8304 14884 8313
rect 15016 8304 15068 8356
rect 16304 8304 16356 8356
rect 17868 8372 17920 8424
rect 18052 8347 18104 8356
rect 9864 8236 9916 8288
rect 12624 8236 12676 8288
rect 12992 8236 13044 8288
rect 13268 8236 13320 8288
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18144 8347 18196 8356
rect 18144 8313 18153 8347
rect 18153 8313 18187 8347
rect 18187 8313 18196 8347
rect 18144 8304 18196 8313
rect 18696 8304 18748 8356
rect 21364 8440 21416 8492
rect 21916 8440 21968 8492
rect 22376 8440 22428 8492
rect 23664 8508 23716 8560
rect 23572 8483 23624 8492
rect 23572 8449 23582 8483
rect 23582 8449 23616 8483
rect 23616 8449 23624 8483
rect 23756 8483 23808 8492
rect 23572 8440 23624 8449
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24768 8508 24820 8560
rect 27252 8576 27304 8628
rect 28172 8576 28224 8628
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 24952 8440 25004 8492
rect 25596 8483 25648 8492
rect 25596 8449 25605 8483
rect 25605 8449 25639 8483
rect 25639 8449 25648 8483
rect 25596 8440 25648 8449
rect 25964 8551 26016 8560
rect 25964 8517 25973 8551
rect 25973 8517 26007 8551
rect 26007 8517 26016 8551
rect 25964 8508 26016 8517
rect 23112 8372 23164 8424
rect 26608 8440 26660 8492
rect 27528 8483 27580 8492
rect 27528 8449 27537 8483
rect 27537 8449 27571 8483
rect 27571 8449 27580 8483
rect 27528 8440 27580 8449
rect 27712 8483 27764 8492
rect 27712 8449 27719 8483
rect 27719 8449 27764 8483
rect 27712 8440 27764 8449
rect 26700 8372 26752 8424
rect 26792 8372 26844 8424
rect 27896 8483 27948 8492
rect 27896 8449 27905 8483
rect 27905 8449 27939 8483
rect 27939 8449 27948 8483
rect 27896 8440 27948 8449
rect 28172 8440 28224 8492
rect 29184 8508 29236 8560
rect 28816 8483 28868 8492
rect 28816 8449 28823 8483
rect 28823 8449 28868 8483
rect 28816 8440 28868 8449
rect 28908 8483 28960 8492
rect 28908 8449 28917 8483
rect 28917 8449 28951 8483
rect 28951 8449 28960 8483
rect 28908 8440 28960 8449
rect 30012 8576 30064 8628
rect 30840 8576 30892 8628
rect 32680 8508 32732 8560
rect 30472 8483 30524 8492
rect 30472 8449 30478 8483
rect 30478 8449 30512 8483
rect 30512 8449 30524 8483
rect 30472 8440 30524 8449
rect 31116 8440 31168 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 31484 8440 31536 8492
rect 22376 8347 22428 8356
rect 22376 8313 22385 8347
rect 22385 8313 22419 8347
rect 22419 8313 22428 8347
rect 22376 8304 22428 8313
rect 22652 8304 22704 8356
rect 22836 8347 22888 8356
rect 22836 8313 22845 8347
rect 22845 8313 22879 8347
rect 22879 8313 22888 8347
rect 22836 8304 22888 8313
rect 30564 8372 30616 8424
rect 30748 8372 30800 8424
rect 33232 8508 33284 8560
rect 33508 8508 33560 8560
rect 33140 8440 33192 8492
rect 24860 8347 24912 8356
rect 24860 8313 24869 8347
rect 24869 8313 24903 8347
rect 24903 8313 24912 8347
rect 24860 8304 24912 8313
rect 25504 8304 25556 8356
rect 27988 8304 28040 8356
rect 28954 8304 29006 8356
rect 29276 8347 29328 8356
rect 29276 8313 29285 8347
rect 29285 8313 29319 8347
rect 29319 8313 29328 8347
rect 29276 8304 29328 8313
rect 29368 8304 29420 8356
rect 33324 8304 33376 8356
rect 33600 8415 33652 8424
rect 33600 8381 33609 8415
rect 33609 8381 33643 8415
rect 33643 8381 33652 8415
rect 34428 8576 34480 8628
rect 34152 8551 34204 8560
rect 34152 8517 34161 8551
rect 34161 8517 34195 8551
rect 34195 8517 34204 8551
rect 34152 8508 34204 8517
rect 34520 8440 34572 8492
rect 34796 8440 34848 8492
rect 35808 8440 35860 8492
rect 33600 8372 33652 8381
rect 35992 8372 36044 8424
rect 17224 8236 17276 8288
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 25596 8236 25648 8288
rect 30012 8236 30064 8288
rect 30380 8236 30432 8288
rect 32312 8236 32364 8288
rect 33416 8236 33468 8288
rect 33968 8304 34020 8356
rect 35624 8304 35676 8356
rect 35532 8279 35584 8288
rect 35532 8245 35541 8279
rect 35541 8245 35575 8279
rect 35575 8245 35584 8279
rect 35532 8236 35584 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 7012 8032 7064 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 7748 7964 7800 8016
rect 8852 8032 8904 8084
rect 5264 7828 5316 7880
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 6184 7871 6236 7880
rect 5356 7828 5408 7837
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 15108 8032 15160 8084
rect 15384 8032 15436 8084
rect 15568 8032 15620 8084
rect 17960 8075 18012 8084
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 18420 8032 18472 8084
rect 18880 8032 18932 8084
rect 23848 8075 23900 8084
rect 23848 8041 23857 8075
rect 23857 8041 23891 8075
rect 23891 8041 23900 8075
rect 23848 8032 23900 8041
rect 24768 8032 24820 8084
rect 25780 8032 25832 8084
rect 26332 8032 26384 8084
rect 26608 8032 26660 8084
rect 28264 8032 28316 8084
rect 28448 8075 28500 8084
rect 28448 8041 28457 8075
rect 28457 8041 28491 8075
rect 28491 8041 28500 8075
rect 28448 8032 28500 8041
rect 28540 8032 28592 8084
rect 30932 8032 30984 8084
rect 31208 8032 31260 8084
rect 31392 8032 31444 8084
rect 35348 8032 35400 8084
rect 7196 7760 7248 7812
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 18604 7896 18656 7948
rect 18696 7896 18748 7948
rect 8484 7692 8536 7744
rect 13176 7760 13228 7812
rect 10048 7692 10100 7744
rect 10508 7692 10560 7744
rect 12440 7692 12492 7744
rect 17868 7760 17920 7812
rect 19064 7828 19116 7880
rect 20996 7871 21048 7880
rect 18052 7760 18104 7812
rect 13360 7692 13412 7744
rect 15108 7692 15160 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 18236 7692 18288 7744
rect 20996 7837 21005 7871
rect 21005 7837 21039 7871
rect 21039 7837 21048 7871
rect 20996 7828 21048 7837
rect 21824 7896 21876 7948
rect 25320 7896 25372 7948
rect 28172 7964 28224 8016
rect 28724 7964 28776 8016
rect 30012 8007 30064 8016
rect 30012 7973 30021 8007
rect 30021 7973 30055 8007
rect 30055 7973 30064 8007
rect 30012 7964 30064 7973
rect 21272 7828 21324 7880
rect 23664 7828 23716 7880
rect 23756 7828 23808 7880
rect 25504 7871 25556 7880
rect 25504 7837 25513 7871
rect 25513 7837 25547 7871
rect 25547 7837 25556 7871
rect 25504 7828 25556 7837
rect 28448 7896 28500 7948
rect 28816 7896 28868 7948
rect 27436 7871 27488 7880
rect 27436 7837 27445 7871
rect 27445 7837 27479 7871
rect 27479 7837 27488 7871
rect 27436 7828 27488 7837
rect 21548 7760 21600 7812
rect 21732 7760 21784 7812
rect 21916 7760 21968 7812
rect 24676 7760 24728 7812
rect 28356 7828 28408 7880
rect 28448 7760 28500 7812
rect 29276 7760 29328 7812
rect 20536 7692 20588 7744
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 21272 7692 21324 7744
rect 23388 7692 23440 7744
rect 24124 7692 24176 7744
rect 27528 7692 27580 7744
rect 28540 7692 28592 7744
rect 32588 7964 32640 8016
rect 30748 7896 30800 7948
rect 30656 7871 30708 7880
rect 30656 7837 30665 7871
rect 30665 7837 30699 7871
rect 30699 7837 30708 7871
rect 30932 7871 30984 7880
rect 30656 7828 30708 7837
rect 30932 7837 30941 7871
rect 30941 7837 30975 7871
rect 30975 7837 30984 7871
rect 30932 7828 30984 7837
rect 31116 7871 31168 7880
rect 31116 7837 31125 7871
rect 31125 7837 31159 7871
rect 31159 7837 31168 7871
rect 31116 7828 31168 7837
rect 31576 7896 31628 7948
rect 32496 7896 32548 7948
rect 34060 7896 34112 7948
rect 32128 7871 32180 7880
rect 32128 7837 32137 7871
rect 32137 7837 32171 7871
rect 32171 7837 32180 7871
rect 32404 7871 32456 7880
rect 32128 7828 32180 7837
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 33232 7828 33284 7880
rect 34612 7828 34664 7880
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 30840 7803 30892 7812
rect 30840 7769 30849 7803
rect 30849 7769 30883 7803
rect 30883 7769 30892 7803
rect 30840 7760 30892 7769
rect 31024 7760 31076 7812
rect 33416 7760 33468 7812
rect 31392 7692 31444 7744
rect 32036 7692 32088 7744
rect 33048 7735 33100 7744
rect 33048 7701 33057 7735
rect 33057 7701 33091 7735
rect 33091 7701 33100 7735
rect 33048 7692 33100 7701
rect 33600 7735 33652 7744
rect 33600 7701 33609 7735
rect 33609 7701 33643 7735
rect 33643 7701 33652 7735
rect 33600 7692 33652 7701
rect 34520 7692 34572 7744
rect 35716 7692 35768 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 6184 7488 6236 7540
rect 8208 7488 8260 7540
rect 9588 7488 9640 7540
rect 5356 7352 5408 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 7748 7395 7800 7404
rect 6000 7284 6052 7336
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 8024 7420 8076 7472
rect 9956 7488 10008 7540
rect 10048 7488 10100 7540
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 7196 7284 7248 7336
rect 9956 7352 10008 7404
rect 10232 7488 10284 7540
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 13544 7488 13596 7497
rect 14464 7488 14516 7540
rect 15108 7488 15160 7540
rect 17960 7488 18012 7540
rect 19064 7488 19116 7540
rect 12624 7420 12676 7472
rect 12532 7352 12584 7404
rect 13452 7352 13504 7404
rect 12716 7284 12768 7336
rect 13268 7284 13320 7336
rect 14924 7352 14976 7404
rect 16396 7420 16448 7472
rect 16764 7420 16816 7472
rect 15384 7352 15436 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 15936 7352 15988 7404
rect 17408 7352 17460 7404
rect 15476 7284 15528 7336
rect 18512 7352 18564 7404
rect 19524 7420 19576 7472
rect 20168 7420 20220 7472
rect 19984 7352 20036 7404
rect 20628 7420 20680 7472
rect 21824 7488 21876 7540
rect 22468 7488 22520 7540
rect 21272 7395 21324 7404
rect 20168 7284 20220 7336
rect 9864 7216 9916 7268
rect 10048 7216 10100 7268
rect 14924 7216 14976 7268
rect 18880 7259 18932 7268
rect 18880 7225 18889 7259
rect 18889 7225 18923 7259
rect 18923 7225 18932 7259
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 24400 7420 24452 7472
rect 22468 7352 22520 7404
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 22008 7284 22060 7336
rect 22744 7284 22796 7336
rect 23388 7352 23440 7404
rect 23940 7352 23992 7404
rect 24860 7488 24912 7540
rect 27344 7488 27396 7540
rect 27896 7488 27948 7540
rect 29000 7488 29052 7540
rect 30748 7488 30800 7540
rect 30932 7488 30984 7540
rect 31392 7488 31444 7540
rect 35348 7488 35400 7540
rect 26792 7420 26844 7472
rect 27436 7420 27488 7472
rect 24860 7352 24912 7404
rect 25596 7395 25648 7404
rect 18880 7216 18932 7225
rect 21456 7216 21508 7268
rect 21916 7259 21968 7268
rect 21916 7225 21925 7259
rect 21925 7225 21959 7259
rect 21959 7225 21968 7259
rect 21916 7216 21968 7225
rect 6552 7148 6604 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 9680 7148 9732 7200
rect 12808 7148 12860 7200
rect 14372 7148 14424 7200
rect 15844 7148 15896 7200
rect 16212 7148 16264 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 20536 7148 20588 7200
rect 23388 7216 23440 7268
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 31852 7420 31904 7472
rect 26056 7284 26108 7336
rect 27068 7327 27120 7336
rect 27068 7293 27077 7327
rect 27077 7293 27111 7327
rect 27111 7293 27120 7327
rect 27068 7284 27120 7293
rect 23572 7216 23624 7268
rect 25596 7148 25648 7200
rect 26792 7216 26844 7268
rect 29828 7395 29880 7404
rect 29828 7361 29837 7395
rect 29837 7361 29871 7395
rect 29871 7361 29880 7395
rect 29828 7352 29880 7361
rect 32312 7352 32364 7404
rect 33048 7420 33100 7472
rect 35532 7420 35584 7472
rect 33600 7352 33652 7404
rect 34704 7395 34756 7404
rect 34704 7361 34713 7395
rect 34713 7361 34747 7395
rect 34747 7361 34756 7395
rect 34704 7352 34756 7361
rect 28632 7148 28684 7200
rect 33968 7191 34020 7200
rect 33968 7157 33977 7191
rect 33977 7157 34011 7191
rect 34011 7157 34020 7191
rect 33968 7148 34020 7157
rect 35900 7148 35952 7200
rect 35992 7148 36044 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5172 6944 5224 6996
rect 6828 6944 6880 6996
rect 13176 6944 13228 6996
rect 17500 6944 17552 6996
rect 10232 6876 10284 6928
rect 12440 6876 12492 6928
rect 16212 6919 16264 6928
rect 4896 6808 4948 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 8208 6808 8260 6860
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 11704 6808 11756 6860
rect 12348 6808 12400 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 7564 6740 7616 6792
rect 8668 6740 8720 6792
rect 6368 6672 6420 6724
rect 7288 6715 7340 6724
rect 7288 6681 7297 6715
rect 7297 6681 7331 6715
rect 7331 6681 7340 6715
rect 7288 6672 7340 6681
rect 8024 6672 8076 6724
rect 9680 6740 9732 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 12716 6740 12768 6792
rect 16212 6885 16221 6919
rect 16221 6885 16255 6919
rect 16255 6885 16264 6919
rect 16212 6876 16264 6885
rect 16396 6876 16448 6928
rect 18420 6944 18472 6996
rect 21180 6944 21232 6996
rect 14280 6808 14332 6860
rect 18052 6851 18104 6860
rect 9404 6672 9456 6724
rect 12256 6672 12308 6724
rect 13820 6740 13872 6792
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 19708 6876 19760 6928
rect 22652 6944 22704 6996
rect 22928 6987 22980 6996
rect 22928 6953 22937 6987
rect 22937 6953 22971 6987
rect 22971 6953 22980 6987
rect 22928 6944 22980 6953
rect 23572 6944 23624 6996
rect 18420 6808 18472 6860
rect 22560 6876 22612 6928
rect 26516 6944 26568 6996
rect 27436 6944 27488 6996
rect 27528 6944 27580 6996
rect 31576 6944 31628 6996
rect 31484 6876 31536 6928
rect 7840 6604 7892 6656
rect 9772 6604 9824 6656
rect 14188 6672 14240 6724
rect 14372 6715 14424 6724
rect 14372 6681 14381 6715
rect 14381 6681 14415 6715
rect 14415 6681 14424 6715
rect 14372 6672 14424 6681
rect 15108 6672 15160 6724
rect 18696 6740 18748 6792
rect 19708 6740 19760 6792
rect 21916 6740 21968 6792
rect 22652 6740 22704 6792
rect 23940 6808 23992 6860
rect 24400 6851 24452 6860
rect 24400 6817 24409 6851
rect 24409 6817 24443 6851
rect 24443 6817 24452 6851
rect 24400 6808 24452 6817
rect 24584 6808 24636 6860
rect 27344 6808 27396 6860
rect 24676 6740 24728 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 25136 6740 25188 6792
rect 25596 6740 25648 6792
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 18236 6715 18288 6724
rect 13728 6604 13780 6656
rect 14648 6604 14700 6656
rect 14832 6604 14884 6656
rect 18236 6681 18245 6715
rect 18245 6681 18279 6715
rect 18279 6681 18288 6715
rect 18236 6672 18288 6681
rect 18328 6715 18380 6724
rect 18328 6681 18337 6715
rect 18337 6681 18371 6715
rect 18371 6681 18380 6715
rect 18328 6672 18380 6681
rect 17868 6604 17920 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 20904 6672 20956 6724
rect 23112 6672 23164 6724
rect 26884 6740 26936 6792
rect 27068 6740 27120 6792
rect 27436 6740 27488 6792
rect 27896 6740 27948 6792
rect 28540 6740 28592 6792
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 30656 6808 30708 6860
rect 31208 6851 31260 6860
rect 31208 6817 31217 6851
rect 31217 6817 31251 6851
rect 31251 6817 31260 6851
rect 31208 6808 31260 6817
rect 31852 6944 31904 6996
rect 32312 6944 32364 6996
rect 32404 6944 32456 6996
rect 35716 6944 35768 6996
rect 35900 6987 35952 6996
rect 35900 6953 35909 6987
rect 35909 6953 35943 6987
rect 35943 6953 35952 6987
rect 35900 6944 35952 6953
rect 30196 6783 30248 6792
rect 30196 6749 30205 6783
rect 30205 6749 30239 6783
rect 30239 6749 30248 6783
rect 30196 6740 30248 6749
rect 30472 6783 30524 6792
rect 30472 6749 30481 6783
rect 30481 6749 30515 6783
rect 30515 6749 30524 6783
rect 30472 6740 30524 6749
rect 33140 6808 33192 6860
rect 35440 6808 35492 6860
rect 27620 6715 27672 6724
rect 27620 6681 27629 6715
rect 27629 6681 27663 6715
rect 27663 6681 27672 6715
rect 27620 6672 27672 6681
rect 27988 6715 28040 6724
rect 27988 6681 27997 6715
rect 27997 6681 28031 6715
rect 28031 6681 28040 6715
rect 27988 6672 28040 6681
rect 28264 6672 28316 6724
rect 33140 6672 33192 6724
rect 33232 6672 33284 6724
rect 34796 6740 34848 6792
rect 35256 6783 35308 6792
rect 35256 6749 35265 6783
rect 35265 6749 35299 6783
rect 35299 6749 35308 6783
rect 35256 6740 35308 6749
rect 36268 6740 36320 6792
rect 36728 6783 36780 6792
rect 36728 6749 36737 6783
rect 36737 6749 36771 6783
rect 36771 6749 36780 6783
rect 36728 6740 36780 6749
rect 37372 6783 37424 6792
rect 37372 6749 37381 6783
rect 37381 6749 37415 6783
rect 37415 6749 37424 6783
rect 37372 6740 37424 6749
rect 35072 6715 35124 6724
rect 35072 6681 35081 6715
rect 35081 6681 35115 6715
rect 35115 6681 35124 6715
rect 35072 6672 35124 6681
rect 35992 6672 36044 6724
rect 22468 6604 22520 6656
rect 22744 6604 22796 6656
rect 24584 6604 24636 6656
rect 28448 6604 28500 6656
rect 30472 6604 30524 6656
rect 30932 6604 30984 6656
rect 31116 6604 31168 6656
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 35900 6604 35952 6656
rect 36268 6604 36320 6656
rect 37188 6647 37240 6656
rect 37188 6613 37197 6647
rect 37197 6613 37231 6647
rect 37231 6613 37240 6647
rect 37188 6604 37240 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4712 6400 4764 6452
rect 6000 6400 6052 6452
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 6460 6400 6512 6452
rect 15568 6400 15620 6452
rect 16028 6443 16080 6452
rect 16028 6409 16037 6443
rect 16037 6409 16071 6443
rect 16071 6409 16080 6443
rect 16028 6400 16080 6409
rect 16672 6400 16724 6452
rect 17224 6400 17276 6452
rect 19248 6400 19300 6452
rect 19984 6400 20036 6452
rect 22468 6400 22520 6452
rect 27160 6400 27212 6452
rect 8392 6332 8444 6384
rect 8944 6375 8996 6384
rect 8944 6341 8953 6375
rect 8953 6341 8987 6375
rect 8987 6341 8996 6375
rect 8944 6332 8996 6341
rect 9220 6332 9272 6384
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7288 6196 7340 6248
rect 8024 6239 8076 6248
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 12532 6332 12584 6384
rect 13544 6332 13596 6384
rect 8208 6264 8260 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 14556 6307 14608 6316
rect 8944 6196 8996 6248
rect 9680 6196 9732 6248
rect 9956 6196 10008 6248
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 14648 6264 14700 6316
rect 14924 6264 14976 6316
rect 16948 6264 17000 6316
rect 20260 6332 20312 6384
rect 21548 6332 21600 6384
rect 22928 6332 22980 6384
rect 17592 6196 17644 6248
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 20628 6196 20680 6248
rect 6920 6128 6972 6180
rect 9036 6128 9088 6180
rect 10140 6128 10192 6180
rect 12532 6128 12584 6180
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 7472 6060 7524 6112
rect 13912 6060 13964 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 16488 6060 16540 6112
rect 18328 6128 18380 6180
rect 20260 6128 20312 6180
rect 21456 6128 21508 6180
rect 22560 6264 22612 6316
rect 24216 6264 24268 6316
rect 26516 6332 26568 6384
rect 27804 6400 27856 6452
rect 29000 6400 29052 6452
rect 27436 6332 27488 6384
rect 26976 6307 27028 6316
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 23572 6128 23624 6180
rect 25136 6196 25188 6248
rect 26976 6273 26985 6307
rect 26985 6273 27019 6307
rect 27019 6273 27028 6307
rect 26976 6264 27028 6273
rect 25228 6128 25280 6180
rect 26516 6196 26568 6248
rect 26792 6196 26844 6248
rect 27344 6307 27396 6316
rect 27344 6273 27353 6307
rect 27353 6273 27387 6307
rect 27387 6273 27396 6307
rect 27344 6264 27396 6273
rect 28080 6264 28132 6316
rect 28264 6307 28316 6316
rect 28264 6273 28273 6307
rect 28273 6273 28307 6307
rect 28307 6273 28316 6307
rect 28264 6264 28316 6273
rect 28540 6264 28592 6316
rect 29644 6332 29696 6384
rect 30196 6400 30248 6452
rect 30288 6332 30340 6384
rect 29368 6307 29420 6316
rect 29368 6273 29402 6307
rect 29402 6273 29420 6307
rect 29368 6264 29420 6273
rect 30380 6264 30432 6316
rect 26700 6128 26752 6180
rect 17500 6060 17552 6112
rect 22652 6060 22704 6112
rect 23388 6060 23440 6112
rect 25964 6060 26016 6112
rect 28448 6128 28500 6180
rect 27436 6060 27488 6112
rect 28356 6060 28408 6112
rect 32036 6332 32088 6384
rect 33048 6332 33100 6384
rect 34796 6400 34848 6452
rect 35164 6400 35216 6452
rect 35624 6400 35676 6452
rect 35072 6332 35124 6384
rect 35808 6400 35860 6452
rect 36268 6332 36320 6384
rect 32680 6264 32732 6316
rect 33140 6307 33192 6316
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 33692 6264 33744 6316
rect 34244 6264 34296 6316
rect 35164 6307 35216 6316
rect 35164 6273 35173 6307
rect 35173 6273 35207 6307
rect 35207 6273 35216 6307
rect 35164 6264 35216 6273
rect 35624 6264 35676 6316
rect 35716 6264 35768 6316
rect 31944 6128 31996 6180
rect 35348 6196 35400 6248
rect 35992 6196 36044 6248
rect 36176 6128 36228 6180
rect 37464 6060 37516 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5632 5856 5684 5908
rect 6460 5788 6512 5840
rect 6920 5788 6972 5840
rect 7564 5788 7616 5840
rect 11888 5856 11940 5908
rect 13728 5856 13780 5908
rect 13820 5856 13872 5908
rect 14924 5899 14976 5908
rect 14924 5865 14933 5899
rect 14933 5865 14967 5899
rect 14967 5865 14976 5899
rect 14924 5856 14976 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 15844 5856 15896 5908
rect 17592 5899 17644 5908
rect 5724 5652 5776 5704
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8760 5652 8812 5704
rect 6736 5584 6788 5636
rect 6828 5584 6880 5636
rect 12164 5652 12216 5704
rect 12716 5652 12768 5704
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 13912 5788 13964 5840
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 16304 5788 16356 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 17316 5788 17368 5840
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 20536 5856 20588 5908
rect 21916 5899 21968 5908
rect 21916 5865 21925 5899
rect 21925 5865 21959 5899
rect 21959 5865 21968 5899
rect 21916 5856 21968 5865
rect 26056 5899 26108 5908
rect 18420 5788 18472 5840
rect 19340 5788 19392 5840
rect 26056 5865 26065 5899
rect 26065 5865 26099 5899
rect 26099 5865 26108 5899
rect 26056 5856 26108 5865
rect 27804 5856 27856 5908
rect 20536 5763 20588 5772
rect 9036 5584 9088 5636
rect 12348 5584 12400 5636
rect 14096 5652 14148 5704
rect 14832 5652 14884 5704
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 14188 5584 14240 5636
rect 15016 5584 15068 5636
rect 17316 5652 17368 5704
rect 20536 5729 20545 5763
rect 20545 5729 20579 5763
rect 20579 5729 20588 5763
rect 20536 5720 20588 5729
rect 18236 5652 18288 5704
rect 18972 5652 19024 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 18328 5584 18380 5636
rect 20168 5652 20220 5704
rect 25964 5788 26016 5840
rect 27620 5788 27672 5840
rect 34244 5856 34296 5908
rect 36176 5856 36228 5908
rect 37832 5788 37884 5840
rect 22560 5763 22612 5772
rect 22560 5729 22569 5763
rect 22569 5729 22603 5763
rect 22603 5729 22612 5763
rect 22560 5720 22612 5729
rect 23020 5720 23072 5772
rect 29828 5763 29880 5772
rect 23664 5652 23716 5704
rect 27252 5652 27304 5704
rect 20628 5584 20680 5636
rect 20904 5584 20956 5636
rect 25688 5584 25740 5636
rect 26240 5584 26292 5636
rect 26884 5584 26936 5636
rect 28080 5652 28132 5704
rect 28540 5695 28592 5704
rect 28540 5661 28549 5695
rect 28549 5661 28583 5695
rect 28583 5661 28592 5695
rect 28540 5652 28592 5661
rect 29828 5729 29837 5763
rect 29837 5729 29871 5763
rect 29871 5729 29880 5763
rect 29828 5720 29880 5729
rect 32128 5720 32180 5772
rect 32588 5720 32640 5772
rect 34704 5763 34756 5772
rect 31024 5652 31076 5704
rect 31760 5652 31812 5704
rect 6460 5516 6512 5568
rect 7104 5516 7156 5568
rect 8024 5516 8076 5568
rect 8300 5516 8352 5568
rect 10232 5516 10284 5568
rect 11796 5516 11848 5568
rect 15108 5516 15160 5568
rect 16304 5516 16356 5568
rect 18604 5559 18656 5568
rect 18604 5525 18613 5559
rect 18613 5525 18647 5559
rect 18647 5525 18656 5559
rect 18604 5516 18656 5525
rect 23112 5516 23164 5568
rect 26516 5516 26568 5568
rect 29000 5584 29052 5636
rect 33416 5652 33468 5704
rect 33692 5695 33744 5704
rect 33692 5661 33701 5695
rect 33701 5661 33735 5695
rect 33735 5661 33744 5695
rect 33692 5652 33744 5661
rect 34704 5729 34713 5763
rect 34713 5729 34747 5763
rect 34747 5729 34756 5763
rect 34704 5720 34756 5729
rect 34612 5652 34664 5704
rect 32680 5627 32732 5636
rect 32680 5593 32689 5627
rect 32689 5593 32723 5627
rect 32723 5593 32732 5627
rect 32680 5584 32732 5593
rect 32864 5627 32916 5636
rect 32864 5593 32873 5627
rect 32873 5593 32907 5627
rect 32907 5593 32916 5627
rect 32864 5584 32916 5593
rect 36728 5671 36780 5704
rect 36728 5652 36737 5671
rect 36737 5652 36771 5671
rect 36771 5652 36780 5671
rect 36084 5584 36136 5636
rect 27804 5516 27856 5568
rect 30840 5516 30892 5568
rect 32588 5516 32640 5568
rect 33876 5516 33928 5568
rect 34244 5516 34296 5568
rect 36912 5516 36964 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 5448 5312 5500 5364
rect 5632 5312 5684 5364
rect 8760 5355 8812 5364
rect 6000 5244 6052 5296
rect 5908 5176 5960 5228
rect 6828 5244 6880 5296
rect 6920 5244 6972 5296
rect 8024 5244 8076 5296
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 6460 5176 6512 5228
rect 7840 5176 7892 5228
rect 9128 5244 9180 5296
rect 9680 5312 9732 5364
rect 6092 5108 6144 5160
rect 8668 5176 8720 5228
rect 10048 5244 10100 5296
rect 10600 5312 10652 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 14556 5312 14608 5364
rect 14924 5312 14976 5364
rect 18328 5312 18380 5364
rect 20536 5312 20588 5364
rect 22468 5312 22520 5364
rect 9496 5185 9501 5212
rect 9501 5185 9535 5212
rect 9535 5185 9548 5212
rect 9496 5160 9548 5185
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 13176 5244 13228 5296
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 12072 5219 12124 5228
rect 11796 5176 11848 5185
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 9128 5108 9180 5160
rect 10784 5108 10836 5160
rect 12808 5176 12860 5228
rect 13820 5176 13872 5228
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 15200 5244 15252 5296
rect 16028 5244 16080 5296
rect 13912 5176 13964 5185
rect 15936 5176 15988 5228
rect 18420 5244 18472 5296
rect 17040 5219 17092 5228
rect 17040 5185 17074 5219
rect 17074 5185 17092 5219
rect 18788 5219 18840 5228
rect 17040 5176 17092 5185
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 19064 5176 19116 5228
rect 20260 5176 20312 5228
rect 23020 5312 23072 5364
rect 23112 5312 23164 5364
rect 26424 5355 26476 5364
rect 26424 5321 26433 5355
rect 26433 5321 26467 5355
rect 26467 5321 26476 5355
rect 26424 5312 26476 5321
rect 22652 5244 22704 5296
rect 20904 5108 20956 5160
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 23296 5219 23348 5228
rect 22284 5176 22336 5185
rect 23296 5185 23305 5219
rect 23305 5185 23339 5219
rect 23339 5185 23348 5219
rect 23296 5176 23348 5185
rect 23480 5176 23532 5228
rect 23848 5176 23900 5228
rect 24124 5176 24176 5228
rect 27436 5312 27488 5364
rect 28264 5312 28316 5364
rect 27620 5244 27672 5296
rect 27712 5244 27764 5296
rect 33232 5312 33284 5364
rect 34244 5355 34296 5364
rect 34244 5321 34253 5355
rect 34253 5321 34287 5355
rect 34287 5321 34296 5355
rect 34244 5312 34296 5321
rect 35624 5312 35676 5364
rect 27252 5219 27304 5228
rect 22192 5108 22244 5160
rect 26424 5108 26476 5160
rect 26884 5108 26936 5160
rect 3516 4972 3568 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 6368 5040 6420 5092
rect 6092 4972 6144 5024
rect 10416 5040 10468 5092
rect 10876 5040 10928 5092
rect 13728 5040 13780 5092
rect 20076 5040 20128 5092
rect 22928 5040 22980 5092
rect 23940 5040 23992 5092
rect 24400 5083 24452 5092
rect 24400 5049 24409 5083
rect 24409 5049 24443 5083
rect 24443 5049 24452 5083
rect 24400 5040 24452 5049
rect 7840 4972 7892 5024
rect 8208 4972 8260 5024
rect 9220 4972 9272 5024
rect 9404 4972 9456 5024
rect 9864 4972 9916 5024
rect 11152 4972 11204 5024
rect 11704 4972 11756 5024
rect 16396 4972 16448 5024
rect 19432 5015 19484 5024
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 20720 4972 20772 5024
rect 25412 4972 25464 5024
rect 26792 4972 26844 5024
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 29276 5219 29328 5228
rect 29276 5185 29285 5219
rect 29285 5185 29319 5219
rect 29319 5185 29328 5219
rect 31300 5244 31352 5296
rect 29276 5176 29328 5185
rect 30656 5176 30708 5228
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 30932 5219 30984 5228
rect 30932 5185 30941 5219
rect 30941 5185 30975 5219
rect 30975 5185 30984 5219
rect 30932 5176 30984 5185
rect 31116 5176 31168 5228
rect 33968 5244 34020 5296
rect 34796 5244 34848 5296
rect 37188 5244 37240 5296
rect 33600 5176 33652 5228
rect 33876 5219 33928 5228
rect 33876 5185 33885 5219
rect 33885 5185 33919 5219
rect 33919 5185 33928 5219
rect 33876 5176 33928 5185
rect 34704 5219 34756 5228
rect 34704 5185 34713 5219
rect 34713 5185 34747 5219
rect 34747 5185 34756 5219
rect 34704 5176 34756 5185
rect 35900 5176 35952 5228
rect 37832 5219 37884 5228
rect 37832 5185 37841 5219
rect 37841 5185 37875 5219
rect 37875 5185 37884 5219
rect 37832 5176 37884 5185
rect 31852 5108 31904 5160
rect 32496 5108 32548 5160
rect 28540 5040 28592 5092
rect 30656 5083 30708 5092
rect 27528 4972 27580 5024
rect 30196 4972 30248 5024
rect 30656 5049 30665 5083
rect 30665 5049 30699 5083
rect 30699 5049 30708 5083
rect 30656 5040 30708 5049
rect 32864 5040 32916 5092
rect 34520 5040 34572 5092
rect 35440 4972 35492 5024
rect 35808 4972 35860 5024
rect 37832 4972 37884 5024
rect 39764 4972 39816 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4988 4768 5040 4820
rect 5448 4700 5500 4752
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 8668 4768 8720 4820
rect 8944 4768 8996 4820
rect 10692 4768 10744 4820
rect 10968 4768 11020 4820
rect 12072 4768 12124 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 12808 4811 12860 4820
rect 12808 4777 12817 4811
rect 12817 4777 12851 4811
rect 12851 4777 12860 4811
rect 12808 4768 12860 4777
rect 12900 4768 12952 4820
rect 14648 4768 14700 4820
rect 17040 4768 17092 4820
rect 18788 4768 18840 4820
rect 20628 4811 20680 4820
rect 10232 4700 10284 4752
rect 10416 4700 10468 4752
rect 13544 4743 13596 4752
rect 6828 4675 6880 4684
rect 1308 4564 1360 4616
rect 4160 4564 4212 4616
rect 5172 4564 5224 4616
rect 6092 4564 6144 4616
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 8300 4632 8352 4684
rect 6920 4564 6972 4616
rect 7104 4607 7156 4616
rect 7104 4573 7138 4607
rect 7138 4573 7156 4607
rect 7104 4564 7156 4573
rect 7380 4564 7432 4616
rect 10600 4632 10652 4684
rect 12992 4632 13044 4684
rect 13544 4709 13553 4743
rect 13553 4709 13587 4743
rect 13587 4709 13596 4743
rect 13544 4700 13596 4709
rect 15936 4700 15988 4752
rect 9864 4564 9916 4616
rect 10324 4564 10376 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 12532 4607 12584 4616
rect 10508 4564 10560 4573
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13176 4564 13228 4616
rect 15568 4632 15620 4684
rect 17040 4632 17092 4684
rect 18328 4632 18380 4684
rect 18420 4632 18472 4684
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 20628 4777 20637 4811
rect 20637 4777 20671 4811
rect 20671 4777 20680 4811
rect 20628 4768 20680 4777
rect 23848 4811 23900 4820
rect 23848 4777 23857 4811
rect 23857 4777 23891 4811
rect 23891 4777 23900 4811
rect 23848 4768 23900 4777
rect 22468 4675 22520 4684
rect 15016 4564 15068 4616
rect 15292 4564 15344 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 5356 4496 5408 4548
rect 10232 4539 10284 4548
rect 1860 4428 1912 4480
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 8760 4428 8812 4480
rect 10232 4505 10241 4539
rect 10241 4505 10275 4539
rect 10275 4505 10284 4539
rect 10232 4496 10284 4505
rect 10968 4496 11020 4548
rect 11152 4539 11204 4548
rect 11152 4505 11161 4539
rect 11161 4505 11195 4539
rect 11195 4505 11204 4539
rect 11152 4496 11204 4505
rect 10784 4428 10836 4480
rect 11060 4428 11112 4480
rect 11612 4496 11664 4548
rect 11796 4496 11848 4548
rect 12716 4496 12768 4548
rect 16488 4496 16540 4548
rect 19064 4564 19116 4616
rect 19984 4564 20036 4616
rect 20812 4564 20864 4616
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 22468 4641 22477 4675
rect 22477 4641 22511 4675
rect 22511 4641 22520 4675
rect 22468 4632 22520 4641
rect 22560 4564 22612 4616
rect 23020 4564 23072 4616
rect 20444 4496 20496 4548
rect 20996 4496 21048 4548
rect 13452 4428 13504 4480
rect 14280 4471 14332 4480
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 19984 4428 20036 4480
rect 20168 4428 20220 4480
rect 21824 4428 21876 4480
rect 23388 4496 23440 4548
rect 23940 4564 23992 4616
rect 26424 4768 26476 4820
rect 26700 4811 26752 4820
rect 26700 4777 26709 4811
rect 26709 4777 26743 4811
rect 26743 4777 26752 4811
rect 26700 4768 26752 4777
rect 26792 4768 26844 4820
rect 28080 4768 28132 4820
rect 29460 4768 29512 4820
rect 29644 4768 29696 4820
rect 31116 4768 31168 4820
rect 33140 4768 33192 4820
rect 33600 4811 33652 4820
rect 33600 4777 33609 4811
rect 33609 4777 33643 4811
rect 33643 4777 33652 4811
rect 33600 4768 33652 4777
rect 37372 4768 37424 4820
rect 37280 4700 37332 4752
rect 27712 4632 27764 4684
rect 28080 4632 28132 4684
rect 25412 4607 25464 4616
rect 25412 4573 25421 4607
rect 25421 4573 25455 4607
rect 25455 4573 25464 4607
rect 25412 4564 25464 4573
rect 24860 4496 24912 4548
rect 27528 4564 27580 4616
rect 28356 4564 28408 4616
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 29000 4564 29052 4616
rect 29828 4632 29880 4684
rect 31484 4607 31536 4616
rect 26056 4539 26108 4548
rect 25136 4428 25188 4480
rect 26056 4505 26065 4539
rect 26065 4505 26099 4539
rect 26099 4505 26108 4539
rect 26056 4496 26108 4505
rect 28264 4496 28316 4548
rect 31484 4573 31493 4607
rect 31493 4573 31527 4607
rect 31527 4573 31536 4607
rect 31484 4564 31536 4573
rect 32220 4607 32272 4616
rect 32220 4573 32229 4607
rect 32229 4573 32263 4607
rect 32263 4573 32272 4607
rect 32220 4564 32272 4573
rect 36912 4632 36964 4684
rect 35716 4564 35768 4616
rect 35808 4607 35860 4616
rect 35808 4573 35817 4607
rect 35817 4573 35851 4607
rect 35851 4573 35860 4607
rect 36452 4607 36504 4616
rect 35808 4564 35860 4573
rect 36452 4573 36461 4607
rect 36461 4573 36495 4607
rect 36495 4573 36504 4607
rect 36452 4564 36504 4573
rect 36544 4564 36596 4616
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 27528 4428 27580 4480
rect 28448 4428 28500 4480
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 29736 4428 29788 4480
rect 30288 4428 30340 4480
rect 31024 4428 31076 4480
rect 31576 4471 31628 4480
rect 31576 4437 31585 4471
rect 31585 4437 31619 4471
rect 31619 4437 31628 4471
rect 31576 4428 31628 4437
rect 33876 4496 33928 4548
rect 36268 4496 36320 4548
rect 32312 4428 32364 4480
rect 35624 4471 35676 4480
rect 35624 4437 35633 4471
rect 35633 4437 35667 4471
rect 35667 4437 35676 4471
rect 35624 4428 35676 4437
rect 37832 4428 37884 4480
rect 39028 4428 39080 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 5632 4267 5684 4276
rect 940 4088 992 4140
rect 3608 4088 3660 4140
rect 5080 4156 5132 4208
rect 5632 4233 5641 4267
rect 5641 4233 5675 4267
rect 5675 4233 5684 4267
rect 5632 4224 5684 4233
rect 7104 4199 7156 4208
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 7104 4165 7113 4199
rect 7113 4165 7147 4199
rect 7147 4165 7156 4199
rect 7104 4156 7156 4165
rect 4528 4088 4580 4097
rect 6736 4088 6788 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7656 4088 7708 4140
rect 4712 4020 4764 4072
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8852 4224 8904 4276
rect 8208 4088 8260 4140
rect 9312 4088 9364 4140
rect 9634 4224 9686 4276
rect 12716 4156 12768 4208
rect 13728 4224 13780 4276
rect 16396 4224 16448 4276
rect 20168 4224 20220 4276
rect 22652 4224 22704 4276
rect 25412 4224 25464 4276
rect 9680 4131 9732 4140
rect 9680 4097 9719 4131
rect 9719 4097 9732 4131
rect 9680 4088 9732 4097
rect 9220 4020 9272 4072
rect 10048 4088 10100 4140
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 12164 4131 12216 4140
rect 10876 4063 10928 4072
rect 2412 3995 2464 4004
rect 2412 3961 2421 3995
rect 2421 3961 2455 3995
rect 2455 3961 2464 3995
rect 2412 3952 2464 3961
rect 2872 3995 2924 4004
rect 2872 3961 2881 3995
rect 2881 3961 2915 3995
rect 2915 3961 2924 3995
rect 2872 3952 2924 3961
rect 3056 3952 3108 4004
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 10048 3952 10100 4004
rect 10600 3952 10652 4004
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 15292 4156 15344 4208
rect 11428 4020 11480 4072
rect 14188 4088 14240 4140
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16764 4088 16816 4140
rect 19064 4156 19116 4208
rect 14280 4020 14332 4072
rect 11152 3952 11204 4004
rect 15108 4020 15160 4072
rect 2044 3884 2096 3936
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 4620 3884 4672 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5816 3884 5868 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 7932 3884 7984 3936
rect 9036 3884 9088 3936
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 12900 3884 12952 3936
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 15016 3952 15068 4004
rect 18880 4088 18932 4140
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 20076 4088 20128 4140
rect 20996 4156 21048 4208
rect 21088 4131 21140 4140
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 21640 4088 21692 4140
rect 21548 4020 21600 4072
rect 22100 4088 22152 4140
rect 22192 4131 22244 4140
rect 22192 4097 22201 4131
rect 22201 4097 22235 4131
rect 22235 4097 22244 4131
rect 25780 4156 25832 4208
rect 22192 4088 22244 4097
rect 23480 4088 23532 4140
rect 23940 4131 23992 4140
rect 23940 4097 23949 4131
rect 23949 4097 23983 4131
rect 23983 4097 23992 4131
rect 23940 4088 23992 4097
rect 24860 4088 24912 4140
rect 26056 4224 26108 4276
rect 27528 4224 27580 4276
rect 28724 4267 28776 4276
rect 28724 4233 28733 4267
rect 28733 4233 28767 4267
rect 28767 4233 28776 4267
rect 28724 4224 28776 4233
rect 29000 4224 29052 4276
rect 28816 4156 28868 4208
rect 29644 4156 29696 4208
rect 25964 4088 26016 4140
rect 26148 4131 26200 4140
rect 26148 4097 26157 4131
rect 26157 4097 26191 4131
rect 26191 4097 26200 4131
rect 26148 4088 26200 4097
rect 26792 4088 26844 4140
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 27804 4131 27856 4140
rect 27804 4097 27813 4131
rect 27813 4097 27847 4131
rect 27847 4097 27856 4131
rect 27804 4088 27856 4097
rect 27988 4131 28040 4140
rect 27988 4097 27997 4131
rect 27997 4097 28031 4131
rect 28031 4097 28040 4131
rect 27988 4088 28040 4097
rect 28264 4088 28316 4140
rect 28908 4131 28960 4140
rect 28908 4097 28917 4131
rect 28917 4097 28951 4131
rect 28951 4097 28960 4131
rect 28908 4088 28960 4097
rect 29092 4088 29144 4140
rect 29276 4131 29328 4140
rect 29276 4097 29285 4131
rect 29285 4097 29319 4131
rect 29319 4097 29328 4131
rect 29276 4088 29328 4097
rect 30748 4088 30800 4140
rect 30840 4131 30892 4140
rect 30840 4097 30849 4131
rect 30849 4097 30883 4131
rect 30883 4097 30892 4131
rect 30840 4088 30892 4097
rect 31300 4088 31352 4140
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 32312 4131 32364 4140
rect 32312 4097 32321 4131
rect 32321 4097 32355 4131
rect 32355 4097 32364 4131
rect 32312 4088 32364 4097
rect 32588 4088 32640 4140
rect 33140 4088 33192 4140
rect 33508 4131 33560 4140
rect 33508 4097 33517 4131
rect 33517 4097 33551 4131
rect 33551 4097 33560 4131
rect 33508 4088 33560 4097
rect 34060 4088 34112 4140
rect 35624 4156 35676 4208
rect 17960 3952 18012 4004
rect 23204 4020 23256 4072
rect 25136 4020 25188 4072
rect 25780 4020 25832 4072
rect 22192 3952 22244 4004
rect 29000 3952 29052 4004
rect 16488 3884 16540 3936
rect 16856 3884 16908 3936
rect 18236 3884 18288 3936
rect 19156 3927 19208 3936
rect 19156 3893 19165 3927
rect 19165 3893 19199 3927
rect 19199 3893 19208 3927
rect 19156 3884 19208 3893
rect 22560 3884 22612 3936
rect 24400 3884 24452 3936
rect 28632 3884 28684 3936
rect 30840 3952 30892 4004
rect 31116 3952 31168 4004
rect 31208 3952 31260 4004
rect 32956 4020 33008 4072
rect 35072 4131 35124 4140
rect 35072 4097 35081 4131
rect 35081 4097 35115 4131
rect 35115 4097 35124 4131
rect 35072 4088 35124 4097
rect 36636 4131 36688 4140
rect 35900 4020 35952 4072
rect 36636 4097 36645 4131
rect 36645 4097 36679 4131
rect 36679 4097 36688 4131
rect 36636 4088 36688 4097
rect 37832 4131 37884 4140
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 29644 3884 29696 3936
rect 31392 3927 31444 3936
rect 31392 3893 31401 3927
rect 31401 3893 31435 3927
rect 31435 3893 31444 3927
rect 31392 3884 31444 3893
rect 32496 3884 32548 3936
rect 32680 3884 32732 3936
rect 33876 3884 33928 3936
rect 34612 3884 34664 3936
rect 35348 3884 35400 3936
rect 38292 3884 38344 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 3148 3680 3200 3732
rect 3056 3655 3108 3664
rect 3056 3621 3065 3655
rect 3065 3621 3099 3655
rect 3099 3621 3108 3655
rect 3056 3612 3108 3621
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 5540 3612 5592 3664
rect 6920 3680 6972 3732
rect 10232 3680 10284 3732
rect 3700 3544 3752 3596
rect 4896 3476 4948 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 4988 3408 5040 3460
rect 5264 3340 5316 3392
rect 6552 3544 6604 3596
rect 6368 3476 6420 3528
rect 6828 3476 6880 3528
rect 5632 3408 5684 3460
rect 7380 3408 7432 3460
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 8668 3544 8720 3596
rect 7656 3476 7708 3485
rect 8300 3476 8352 3528
rect 8852 3544 8904 3596
rect 10232 3544 10284 3596
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9036 3476 9088 3528
rect 9496 3476 9548 3528
rect 11152 3544 11204 3596
rect 12624 3680 12676 3732
rect 14740 3680 14792 3732
rect 16120 3680 16172 3732
rect 21548 3723 21600 3732
rect 21548 3689 21557 3723
rect 21557 3689 21591 3723
rect 21591 3689 21600 3723
rect 21548 3680 21600 3689
rect 12716 3612 12768 3664
rect 13820 3544 13872 3596
rect 19248 3587 19300 3596
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 22468 3680 22520 3732
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 26332 3680 26384 3732
rect 26792 3723 26844 3732
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 23204 3544 23256 3596
rect 28264 3680 28316 3732
rect 29276 3680 29328 3732
rect 29368 3680 29420 3732
rect 28816 3612 28868 3664
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 12164 3476 12216 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 15200 3476 15252 3528
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16488 3476 16540 3528
rect 8208 3408 8260 3460
rect 11152 3408 11204 3460
rect 11980 3408 12032 3460
rect 15752 3408 15804 3460
rect 16764 3408 16816 3460
rect 17316 3408 17368 3460
rect 19340 3476 19392 3528
rect 20996 3408 21048 3460
rect 21732 3476 21784 3528
rect 22836 3476 22888 3528
rect 24952 3476 25004 3528
rect 27528 3476 27580 3528
rect 22192 3408 22244 3460
rect 25228 3408 25280 3460
rect 27344 3408 27396 3460
rect 28724 3544 28776 3596
rect 29276 3544 29328 3596
rect 28172 3476 28224 3528
rect 33508 3680 33560 3732
rect 33876 3680 33928 3732
rect 34704 3680 34756 3732
rect 36452 3680 36504 3732
rect 36636 3612 36688 3664
rect 32312 3544 32364 3596
rect 32956 3587 33008 3596
rect 27988 3408 28040 3460
rect 29184 3408 29236 3460
rect 32220 3476 32272 3528
rect 32404 3476 32456 3528
rect 32956 3553 32965 3587
rect 32965 3553 32999 3587
rect 32999 3553 33008 3587
rect 32956 3544 33008 3553
rect 33048 3544 33100 3596
rect 33140 3519 33192 3528
rect 30656 3408 30708 3460
rect 31392 3408 31444 3460
rect 31484 3408 31536 3460
rect 7656 3340 7708 3392
rect 7840 3340 7892 3392
rect 10508 3340 10560 3392
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 24860 3340 24912 3392
rect 30840 3340 30892 3392
rect 32312 3408 32364 3460
rect 33140 3485 33149 3519
rect 33149 3485 33183 3519
rect 33183 3485 33192 3519
rect 33140 3476 33192 3485
rect 34980 3544 35032 3596
rect 35624 3544 35676 3596
rect 34796 3476 34848 3528
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 36176 3476 36228 3528
rect 32588 3340 32640 3392
rect 33232 3408 33284 3460
rect 34520 3340 34572 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 36084 3340 36136 3392
rect 37556 3340 37608 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2688 3136 2740 3188
rect 3240 3136 3292 3188
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 4436 3000 4488 3052
rect 5448 3068 5500 3120
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 6552 3136 6604 3188
rect 7840 3136 7892 3188
rect 8024 3136 8076 3188
rect 10324 3136 10376 3188
rect 10692 3136 10744 3188
rect 11152 3136 11204 3188
rect 13636 3136 13688 3188
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 6644 3111 6696 3120
rect 6644 3077 6678 3111
rect 6678 3077 6696 3111
rect 6644 3068 6696 3077
rect 5540 3000 5592 3052
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 4620 2932 4672 2984
rect 7196 3000 7248 3052
rect 8300 3000 8352 3052
rect 8944 3068 8996 3120
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9680 3000 9732 3052
rect 10232 3000 10284 3052
rect 12164 3068 12216 3120
rect 13912 3111 13964 3120
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 12072 3043 12124 3052
rect 12072 3009 12106 3043
rect 12106 3009 12124 3043
rect 12072 3000 12124 3009
rect 13176 3000 13228 3052
rect 13728 3000 13780 3052
rect 14924 3111 14976 3120
rect 14924 3077 14933 3111
rect 14933 3077 14967 3111
rect 14967 3077 14976 3111
rect 14924 3068 14976 3077
rect 14740 3000 14792 3052
rect 16672 3136 16724 3188
rect 20444 3136 20496 3188
rect 20904 3136 20956 3188
rect 15292 3000 15344 3052
rect 2228 2907 2280 2916
rect 2228 2873 2237 2907
rect 2237 2873 2271 2907
rect 2271 2873 2280 2907
rect 2228 2864 2280 2873
rect 7656 2864 7708 2916
rect 15108 2932 15160 2984
rect 8668 2907 8720 2916
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 4068 2796 4120 2848
rect 5080 2796 5132 2848
rect 8668 2873 8677 2907
rect 8677 2873 8711 2907
rect 8711 2873 8720 2907
rect 8668 2864 8720 2873
rect 9588 2864 9640 2916
rect 7932 2796 7984 2848
rect 8944 2796 8996 2848
rect 10600 2796 10652 2848
rect 11980 2796 12032 2848
rect 14096 2864 14148 2916
rect 16764 3068 16816 3120
rect 17224 3068 17276 3120
rect 19064 3068 19116 3120
rect 23572 3136 23624 3188
rect 25780 3136 25832 3188
rect 27804 3136 27856 3188
rect 30472 3136 30524 3188
rect 16396 3000 16448 3052
rect 19156 3000 19208 3052
rect 20628 3000 20680 3052
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 22376 3000 22428 3052
rect 20352 2932 20404 2984
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 23204 3043 23256 3052
rect 23204 3009 23213 3043
rect 23213 3009 23247 3043
rect 23247 3009 23256 3043
rect 23204 3000 23256 3009
rect 23296 3043 23348 3052
rect 23296 3009 23305 3043
rect 23305 3009 23339 3043
rect 23339 3009 23348 3043
rect 23296 3000 23348 3009
rect 24584 3000 24636 3052
rect 24860 3043 24912 3052
rect 24860 3009 24869 3043
rect 24869 3009 24903 3043
rect 24903 3009 24912 3043
rect 24860 3000 24912 3009
rect 21824 2932 21876 2941
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 13820 2796 13872 2848
rect 14280 2796 14332 2848
rect 28172 3068 28224 3120
rect 25964 3000 26016 3052
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 26516 2932 26568 2984
rect 27712 3000 27764 3052
rect 27896 3000 27948 3052
rect 28356 3000 28408 3052
rect 27988 2932 28040 2984
rect 28816 2932 28868 2984
rect 32496 3136 32548 3188
rect 34520 3136 34572 3188
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 30932 3000 30984 3052
rect 31116 3043 31168 3052
rect 31116 3009 31125 3043
rect 31125 3009 31159 3043
rect 31159 3009 31168 3043
rect 31116 3000 31168 3009
rect 31300 3000 31352 3052
rect 32404 3043 32456 3052
rect 32404 3009 32413 3043
rect 32413 3009 32447 3043
rect 32447 3009 32456 3043
rect 32404 3000 32456 3009
rect 32680 3043 32732 3052
rect 32680 3009 32714 3043
rect 32714 3009 32732 3043
rect 32680 3000 32732 3009
rect 29828 2932 29880 2984
rect 31208 2975 31260 2984
rect 31208 2941 31217 2975
rect 31217 2941 31251 2975
rect 31251 2941 31260 2975
rect 31208 2932 31260 2941
rect 33784 2932 33836 2984
rect 36360 3136 36412 3188
rect 34796 3068 34848 3120
rect 34980 3043 35032 3052
rect 34980 3009 34989 3043
rect 34989 3009 35023 3043
rect 35023 3009 35032 3043
rect 34980 3000 35032 3009
rect 35808 3068 35860 3120
rect 35440 2932 35492 2984
rect 35992 3000 36044 3052
rect 36636 3000 36688 3052
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 36544 2932 36596 2984
rect 37464 2932 37516 2984
rect 27068 2864 27120 2916
rect 29000 2864 29052 2916
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 18144 2796 18196 2848
rect 21824 2796 21876 2848
rect 23112 2796 23164 2848
rect 24860 2796 24912 2848
rect 25228 2796 25280 2848
rect 28172 2796 28224 2848
rect 28540 2796 28592 2848
rect 29276 2796 29328 2848
rect 33416 2864 33468 2916
rect 34796 2864 34848 2916
rect 32772 2796 32824 2848
rect 33140 2796 33192 2848
rect 36176 2796 36228 2848
rect 36820 2796 36872 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6644 2592 6696 2644
rect 7380 2592 7432 2644
rect 8116 2635 8168 2644
rect 2136 2524 2188 2576
rect 4712 2524 4764 2576
rect 5172 2524 5224 2576
rect 7472 2524 7524 2576
rect 6920 2456 6972 2508
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 9312 2635 9364 2644
rect 9312 2601 9321 2635
rect 9321 2601 9355 2635
rect 9355 2601 9364 2635
rect 9312 2592 9364 2601
rect 10968 2592 11020 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 15844 2635 15896 2644
rect 15844 2601 15853 2635
rect 15853 2601 15887 2635
rect 15887 2601 15896 2635
rect 15844 2592 15896 2601
rect 18696 2592 18748 2644
rect 22192 2592 22244 2644
rect 28080 2592 28132 2644
rect 28356 2592 28408 2644
rect 17316 2524 17368 2576
rect 17408 2524 17460 2576
rect 21088 2524 21140 2576
rect 25596 2524 25648 2576
rect 29000 2592 29052 2644
rect 30472 2635 30524 2644
rect 30472 2601 30481 2635
rect 30481 2601 30515 2635
rect 30515 2601 30524 2635
rect 30472 2592 30524 2601
rect 29276 2524 29328 2576
rect 29368 2524 29420 2576
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 3884 2388 3936 2440
rect 572 2320 624 2372
rect 4252 2320 4304 2372
rect 8024 2388 8076 2440
rect 9404 2388 9456 2440
rect 10416 2388 10468 2440
rect 10968 2388 11020 2440
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 3148 2252 3200 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 7104 2320 7156 2372
rect 7932 2252 7984 2304
rect 14004 2456 14056 2508
rect 17776 2456 17828 2508
rect 25504 2456 25556 2508
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 15292 2388 15344 2440
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17960 2388 18012 2440
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 19432 2388 19484 2440
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 25044 2388 25096 2440
rect 25136 2388 25188 2440
rect 28448 2456 28500 2508
rect 29644 2456 29696 2508
rect 30104 2456 30156 2508
rect 34520 2592 34572 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 31668 2524 31720 2576
rect 32772 2456 32824 2508
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 30196 2388 30248 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 31576 2388 31628 2440
rect 33416 2388 33468 2440
rect 34612 2456 34664 2508
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 37372 2388 37424 2440
rect 13820 2320 13872 2372
rect 16580 2320 16632 2372
rect 22652 2320 22704 2372
rect 28632 2320 28684 2372
rect 18880 2252 18932 2304
rect 19984 2252 20036 2304
rect 20352 2252 20404 2304
rect 24124 2252 24176 2304
rect 26332 2252 26384 2304
rect 30840 2252 30892 2304
rect 33140 2252 33192 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 5540 2048 5592 2100
rect 8392 2048 8444 2100
rect 9220 2048 9272 2100
rect 14372 2048 14424 2100
rect 2688 1980 2740 2032
rect 12164 1980 12216 2032
rect 2504 1912 2556 1964
rect 3792 1912 3844 1964
rect 18604 2048 18656 2100
rect 11428 1844 11480 1896
rect 6092 1776 6144 1828
rect 9496 1776 9548 1828
rect 5172 1708 5224 1760
rect 11244 1708 11296 1760
rect 204 1640 256 1692
rect 8484 1640 8536 1692
rect 5448 1572 5500 1624
rect 8760 1572 8812 1624
rect 3608 1368 3660 1420
rect 5356 1368 5408 1420
rect 6000 1368 6052 1420
rect 6552 1368 6604 1420
rect 6736 1368 6788 1420
rect 9128 1368 9180 1420
rect 1952 1096 2004 1148
rect 6184 1096 6236 1148
rect 10324 1096 10376 1148
rect 11796 1096 11848 1148
<< metal2 >>
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 23492 16658 23612 16674
rect 23492 16652 23624 16658
rect 23492 16646 23572 16652
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 22664 16114 22692 16390
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 20732 15502 20760 15982
rect 23032 15706 23060 16526
rect 23492 15978 23520 16646
rect 23572 16594 23624 16600
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 28816 16584 28868 16590
rect 28816 16526 28868 16532
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23584 16250 23612 16458
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 20456 14618 20484 14962
rect 20732 14822 20760 15438
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 15162 21864 15370
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21928 14958 21956 15302
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 9508 12306 9536 12582
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11762 5856 12038
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5644 10810 5672 11018
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 204 1692 256 1698
rect 204 1634 256 1640
rect 216 800 244 1634
rect 584 800 612 2314
rect 952 800 980 4082
rect 1320 800 1348 4558
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 3126 1900 4422
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1964 1154 1992 3470
rect 2056 2854 2084 3878
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2148 2582 2176 9590
rect 2240 3738 2268 9658
rect 2424 4010 2452 10542
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 4010 2912 10406
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3146 4448 3202 4457
rect 3068 4010 3096 4422
rect 3146 4383 3202 4392
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3160 3738 3188 4383
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3664 3108 3670
rect 3054 3632 3056 3641
rect 3108 3632 3110 3641
rect 3054 3567 3110 3576
rect 2686 3496 2742 3505
rect 2686 3431 2742 3440
rect 2700 3194 2728 3431
rect 3252 3194 3280 10474
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4080 9178 4108 9590
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4632 8634 4660 8842
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4724 6458 4752 10134
rect 6564 10062 6592 10950
rect 6748 10674 6776 11494
rect 6932 10810 6960 12174
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 7024 11218 7052 11766
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4908 8974 4936 9590
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 6866 4936 8910
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 5092 5914 5120 8366
rect 5368 8294 5396 9930
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5276 7886 5304 8230
rect 5368 7886 5396 8230
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 7410 5396 7822
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2226 2952 2282 2961
rect 2226 2887 2228 2896
rect 2280 2887 2282 2896
rect 2228 2858 2280 2864
rect 2136 2576 2188 2582
rect 2136 2518 2188 2524
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 1970 2544 2246
rect 2700 2038 2728 2382
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 2688 2032 2740 2038
rect 2688 1974 2740 1980
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 1952 1148 2004 1154
rect 1952 1090 2004 1096
rect 3160 800 3188 2246
rect 3528 800 3556 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 5000 4826 5028 4966
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5184 4706 5212 6938
rect 5460 5370 5488 8842
rect 5644 8634 5672 9522
rect 5736 9178 5764 9522
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 8498 5764 9114
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 8090 5580 8298
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5914 5672 6054
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5538 5264 5594 5273
rect 5538 5199 5594 5208
rect 5000 4678 5212 4706
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 1426 3648 4082
rect 4172 3992 4200 4558
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4528 4140 4580 4146
rect 4632 4134 4844 4162
rect 4632 4128 4660 4134
rect 4580 4100 4660 4128
rect 4528 4082 4580 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4080 3964 4200 3992
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3602 3740 3878
rect 4080 3720 4108 3964
rect 4620 3936 4672 3942
rect 4618 3904 4620 3913
rect 4672 3904 4674 3913
rect 4214 3836 4522 3856
rect 4618 3839 4674 3848
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4080 3692 4200 3720
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 4172 3233 4200 3692
rect 4158 3224 4214 3233
rect 4158 3159 4214 3168
rect 4434 3088 4490 3097
rect 4434 3023 4436 3032
rect 4488 3023 4490 3032
rect 4436 2994 4488 3000
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3884 2440 3936 2446
rect 4080 2417 4108 2790
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3884 2382 3936 2388
rect 4066 2408 4122 2417
rect 3804 1970 3832 2382
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3896 800 3924 2382
rect 4066 2343 4122 2352
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4264 800 4292 2314
rect 4632 800 4660 2926
rect 4724 2582 4752 4014
rect 4816 3505 4844 4134
rect 4908 4049 4936 4422
rect 4894 4040 4950 4049
rect 4894 3975 4950 3984
rect 5000 3942 5028 4678
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5354 4584 5410 4593
rect 5078 4312 5134 4321
rect 5078 4247 5134 4256
rect 5092 4214 5120 4247
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4896 3528 4948 3534
rect 4802 3496 4858 3505
rect 4896 3470 4948 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4802 3431 4858 3440
rect 4908 3369 4936 3470
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4894 3360 4950 3369
rect 4894 3295 4950 3304
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 5000 800 5028 3402
rect 5092 2854 5120 3470
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5184 2582 5212 4558
rect 5354 4519 5356 4528
rect 5408 4519 5410 4528
rect 5356 4490 5408 4496
rect 5262 4176 5318 4185
rect 5262 4111 5318 4120
rect 5276 3398 5304 4111
rect 5460 3641 5488 4694
rect 5552 3670 5580 5199
rect 5644 4282 5672 5306
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 3664 5592 3670
rect 5446 3632 5502 3641
rect 5540 3606 5592 3612
rect 5446 3567 5502 3576
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5644 3194 5672 3402
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 1766 5212 2246
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5460 1630 5488 3062
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5552 2106 5580 2994
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5448 1624 5500 1630
rect 5448 1566 5500 1572
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 5368 800 5396 1362
rect 5736 800 5764 5646
rect 5828 4457 5856 9930
rect 6196 9178 6224 9998
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 8566 6316 8910
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6380 8498 6408 9862
rect 6564 9586 6592 9998
rect 6748 9586 6776 10610
rect 6932 9926 6960 10610
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 7024 9654 7052 11154
rect 7668 11150 7696 12038
rect 8312 11694 8340 12242
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11898 8616 12174
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 9232 11762 9260 12038
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7208 10198 7236 10610
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7208 10062 7236 10134
rect 7760 10062 7788 11290
rect 8312 10810 8340 11630
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7944 10266 7972 10610
rect 8312 10606 8340 10746
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8404 10266 8432 11698
rect 9692 11218 9720 12786
rect 10520 12442 10548 12786
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8974 6500 9318
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6656 8362 6684 8978
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7546 6224 7822
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6748 7410 6776 8502
rect 6840 7410 6868 8842
rect 7024 8498 7052 9590
rect 7760 9042 7788 9998
rect 8772 9926 8800 10610
rect 9324 10062 9352 10610
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9466 7880 9522
rect 8392 9512 8444 9518
rect 7852 9438 7972 9466
rect 8392 9454 8444 9460
rect 7944 9382 7972 9438
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 8090 7052 8434
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7208 7818 7236 8774
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 6458 6040 7278
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6380 6458 6408 6666
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 5846 6500 6394
rect 6564 6322 6592 7142
rect 6840 7002 6868 7346
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6932 5846 6960 6122
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3058 5856 3878
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5920 2281 5948 5170
rect 5906 2272 5962 2281
rect 5906 2207 5962 2216
rect 6012 1426 6040 5238
rect 6472 5234 6500 5510
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 5030 6132 5102
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6274 4720 6330 4729
rect 6274 4655 6330 4664
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 1834 6132 4558
rect 6288 3777 6316 4655
rect 6274 3768 6330 3777
rect 6380 3754 6408 5034
rect 6748 4865 6776 5578
rect 6840 5302 6868 5578
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6734 4856 6790 4865
rect 6734 4791 6790 4800
rect 6840 4690 6868 5238
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6458 3768 6514 3777
rect 6380 3726 6458 3754
rect 6274 3703 6330 3712
rect 6458 3703 6514 3712
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6380 3058 6408 3470
rect 6564 3194 6592 3538
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6656 2650 6684 3062
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6748 1426 6776 4082
rect 6840 3534 6868 4626
rect 6932 4622 6960 5238
rect 7116 4622 7144 5510
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6932 3738 6960 4082
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6552 1420 6604 1426
rect 6552 1362 6604 1368
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6184 1148 6236 1154
rect 6184 1090 6236 1096
rect 6196 800 6224 1090
rect 6564 800 6592 1362
rect 6932 800 6960 2450
rect 7116 2378 7144 4150
rect 7208 3058 7236 7278
rect 7300 6730 7328 8230
rect 7484 6866 7512 8910
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7760 7410 7788 7958
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7576 6798 7604 7142
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7852 6662 7880 8434
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7300 800 7328 6190
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5710 7512 6054
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4185 7420 4558
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 2650 7420 3402
rect 7470 2816 7526 2825
rect 7470 2751 7526 2760
rect 7576 2774 7604 5782
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7852 5030 7880 5170
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3534 7696 4082
rect 7852 4078 7880 4966
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7944 3942 7972 9318
rect 8404 9178 8432 9454
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8036 8090 8064 9114
rect 8772 9042 8800 9862
rect 9324 9586 9352 9998
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 9110 9076 9318
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7478 8064 8026
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8036 6254 8064 6666
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5710 8064 6190
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 5574 8064 5646
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3398 7696 3470
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7760 3176 7788 3878
rect 7840 3392 7892 3398
rect 7838 3360 7840 3369
rect 7892 3360 7894 3369
rect 7838 3295 7894 3304
rect 8036 3194 8064 5238
rect 7840 3188 7892 3194
rect 7668 3148 7840 3176
rect 7668 2922 7696 3148
rect 7840 3130 7892 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2582 7512 2751
rect 7576 2746 7696 2774
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7668 800 7696 2746
rect 7944 2310 7972 2790
rect 8128 2650 8156 7346
rect 8220 6866 8248 7482
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 5030 8248 6258
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8220 4146 8248 4762
rect 8312 4690 8340 5510
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 2825 8248 3402
rect 8312 3058 8340 3470
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8206 2816 8262 2825
rect 8206 2751 8262 2760
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8404 2553 8432 6326
rect 8390 2544 8446 2553
rect 8390 2479 8446 2488
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8036 800 8064 2382
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8404 800 8432 2042
rect 8496 1698 8524 7686
rect 8588 7410 8616 8910
rect 8956 8634 8984 8910
rect 9232 8634 9260 8910
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8680 6798 8708 8298
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8772 5370 8800 5646
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8680 4826 8708 5170
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8680 2922 8708 3538
rect 8772 3058 8800 4422
rect 8864 4282 8892 8026
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8956 6390 8984 7511
rect 9232 6390 9260 8570
rect 9416 8498 9444 11086
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9600 10606 9628 10746
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 9994 9536 10406
rect 9784 10266 9812 12174
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 9968 10810 9996 12106
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11830 10456 12038
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10336 10742 10364 11494
rect 10428 11218 10456 11766
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10520 11121 10548 12106
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10506 11112 10562 11121
rect 10704 11082 10732 12038
rect 10506 11047 10562 11056
rect 10692 11076 10744 11082
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 10520 10198 10548 11047
rect 10692 11018 10744 11024
rect 11348 10810 11376 12174
rect 11624 11830 11652 12582
rect 14936 12434 14964 13262
rect 14752 12406 14964 12434
rect 16396 12436 16448 12442
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11440 10674 11468 10950
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9416 6730 9444 8434
rect 9600 7546 9628 8434
rect 9692 7698 9720 9454
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8566 9812 8774
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9692 7670 9812 7698
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6798 9720 7142
rect 9784 6866 9812 7670
rect 9876 7274 9904 8230
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7546 10088 7686
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9968 7410 9996 7482
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9784 6662 9812 6802
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 8956 4826 8984 6190
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9048 5642 9076 6122
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9692 5370 9720 6190
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9128 5296 9180 5302
rect 9494 5264 9550 5273
rect 9128 5238 9180 5244
rect 9140 5166 9168 5238
rect 9477 5208 9494 5250
rect 9477 5188 9496 5208
rect 9128 5160 9180 5166
rect 9548 5199 9550 5208
rect 9496 5154 9548 5160
rect 9180 5120 9444 5148
rect 9128 5102 9180 5108
rect 9416 5114 9444 5120
rect 9692 5114 9720 5306
rect 9876 5137 9904 7210
rect 9968 6254 9996 7346
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10060 6798 10088 7210
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10060 5302 10088 6734
rect 10152 6186 10180 9930
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10428 9178 10456 9522
rect 10612 9178 10640 10610
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10428 8650 10456 9114
rect 10980 8838 11008 9998
rect 11072 9042 11100 10202
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9722 11376 9998
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10428 8622 10548 8650
rect 10520 8566 10548 8622
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10244 6934 10272 7482
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10244 5234 10272 5510
rect 10232 5228 10284 5234
rect 10284 5188 10364 5216
rect 10232 5170 10284 5176
rect 9416 5086 9720 5114
rect 9862 5128 9918 5137
rect 9862 5063 9918 5072
rect 10230 5128 10286 5137
rect 10230 5063 10286 5072
rect 9220 5024 9272 5030
rect 9404 5024 9456 5030
rect 9272 4984 9404 5012
rect 9220 4966 9272 4972
rect 9404 4966 9456 4972
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9876 4622 9904 4966
rect 10244 4758 10272 5063
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10336 4622 10364 5188
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10428 4758 10456 5034
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10520 4622 10548 7686
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10612 4690 10640 5306
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 9864 4616 9916 4622
rect 10324 4616 10376 4622
rect 9864 4558 9916 4564
rect 10138 4584 10194 4593
rect 10324 4558 10376 4564
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10138 4519 10194 4528
rect 10232 4548 10284 4554
rect 9646 4406 10088 4434
rect 9646 4282 9674 4406
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 9634 4276 9686 4282
rect 9634 4218 9686 4224
rect 8864 3602 8892 4218
rect 9678 4176 9734 4185
rect 9312 4140 9364 4146
rect 10060 4146 10088 4406
rect 9678 4111 9680 4120
rect 9312 4082 9364 4088
rect 9732 4111 9734 4120
rect 10048 4140 10100 4146
rect 9680 4082 9732 4088
rect 10048 4082 10100 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 9048 3534 9076 3878
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8956 3126 8984 3470
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8956 2417 8984 2790
rect 8942 2408 8998 2417
rect 8942 2343 8998 2352
rect 9232 2106 9260 4014
rect 9324 2650 9352 4082
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9416 2446 9444 3878
rect 10060 3641 10088 3946
rect 9494 3632 9550 3641
rect 9494 3567 9550 3576
rect 9770 3632 9826 3641
rect 9770 3567 9826 3576
rect 10046 3632 10102 3641
rect 10046 3567 10102 3576
rect 9508 3534 9536 3567
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9784 3176 9812 3567
rect 9600 3148 9812 3176
rect 9600 2922 9628 3148
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9692 2774 9720 2994
rect 10152 2774 10180 4519
rect 10232 4490 10284 4496
rect 10244 4185 10272 4490
rect 10230 4176 10286 4185
rect 10704 4146 10732 4762
rect 10796 4486 10824 5102
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10230 4111 10286 4120
rect 10692 4140 10744 4146
rect 10244 3738 10272 4111
rect 10692 4082 10744 4088
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3058 10272 3538
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9692 2746 9904 2774
rect 10152 2746 10272 2774
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 8484 1692 8536 1698
rect 8484 1634 8536 1640
rect 8760 1624 8812 1630
rect 8760 1566 8812 1572
rect 8772 800 8800 1566
rect 9128 1420 9180 1426
rect 9128 1362 9180 1368
rect 9140 800 9168 1362
rect 9508 800 9536 1770
rect 9876 800 9904 2746
rect 10244 800 10272 2746
rect 10336 1154 10364 3130
rect 10428 2446 10456 3878
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10520 1442 10548 3334
rect 10612 2854 10640 3946
rect 10704 3194 10732 4082
rect 10888 4078 10916 5034
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10980 4554 11008 4762
rect 11164 4554 11192 4966
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10690 3088 10746 3097
rect 10690 3023 10746 3032
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10520 1414 10640 1442
rect 10324 1148 10376 1154
rect 10324 1090 10376 1096
rect 10612 800 10640 1414
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10704 762 10732 3023
rect 10980 2650 11008 3470
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10968 2440 11020 2446
rect 11072 2428 11100 4422
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11164 3602 11192 3946
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3194 11192 3402
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11020 2400 11100 2428
rect 10968 2382 11020 2388
rect 11256 1766 11284 8910
rect 11348 8430 11376 8978
rect 11440 8906 11468 10610
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11532 8974 11560 9862
rect 11624 9722 11652 9862
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9586 11652 9658
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11808 8974 11836 9454
rect 11992 9382 12020 9998
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 8974 12020 9318
rect 12084 9178 12112 12174
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 11014 12388 11698
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10674 12388 10950
rect 12452 10742 12480 12038
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12544 11354 12572 11834
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13280 11558 13308 11766
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12348 10668 12400 10674
rect 12636 10656 12664 11154
rect 12728 10742 12756 11290
rect 13280 11218 13308 11494
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13174 11112 13230 11121
rect 13174 11047 13176 11056
rect 13228 11047 13230 11056
rect 13176 11018 13228 11024
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12348 10610 12400 10616
rect 12544 10628 12664 10656
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12176 9382 12204 10202
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 12544 8838 12572 10628
rect 13280 10062 13308 11154
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13372 9042 13400 11698
rect 13556 9586 13584 11698
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 9178 13584 9522
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12084 8498 12112 8774
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 12360 6866 12388 8774
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 7834 12664 8230
rect 12636 7806 12848 7834
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 6934 12480 7686
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11624 4554 11652 6734
rect 11716 5030 11744 6802
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11900 5914 11928 6258
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11808 4554 11836 5170
rect 12084 4826 12112 5170
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11334 4312 11390 4321
rect 11334 4247 11390 4256
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 10888 870 11008 898
rect 10888 762 10916 870
rect 10980 800 11008 870
rect 11348 800 11376 4247
rect 12176 4146 12204 5646
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 1902 11468 4014
rect 12176 3534 12204 4082
rect 12268 3913 12296 6666
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12254 3904 12310 3913
rect 12254 3839 12310 3848
rect 12164 3528 12216 3534
rect 12360 3516 12388 5578
rect 12452 4826 12480 6870
rect 12544 6390 12572 7346
rect 12636 6866 12664 7414
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12728 6798 12756 7278
rect 12820 7206 12848 7806
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4706 12572 6122
rect 12728 5710 12756 6190
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12912 5370 12940 8842
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12820 4826 12848 5170
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12544 4678 12756 4706
rect 12532 4616 12584 4622
rect 12584 4576 12664 4604
rect 12532 4558 12584 4564
rect 12636 4146 12664 4576
rect 12728 4554 12756 4678
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12716 4208 12768 4214
rect 12912 4196 12940 4762
rect 13004 4690 13032 8230
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7002 13216 7754
rect 13280 7342 13308 8230
rect 13372 7750 13400 8434
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13556 7546 13584 8366
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13464 7290 13492 7346
rect 13740 7290 13768 8502
rect 13832 8362 13860 12174
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14016 11354 14044 11698
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14016 10742 14044 11290
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14200 10062 14228 11494
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 10674 14412 11086
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14292 9994 14320 10542
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14476 9586 14504 11494
rect 14568 10062 14596 11698
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14660 9586 14688 10950
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13280 6882 13308 7278
rect 13464 7262 13768 7290
rect 13188 6854 13308 6882
rect 13188 5710 13216 6854
rect 13740 6662 13768 7262
rect 14292 6866 14320 8910
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14476 7546 14504 8434
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14752 7426 14780 12406
rect 16396 12378 16448 12384
rect 16210 12336 16266 12345
rect 16210 12271 16266 12280
rect 16224 12238 16252 12271
rect 16212 12232 16264 12238
rect 14830 12200 14886 12209
rect 16212 12174 16264 12180
rect 14830 12135 14832 12144
rect 14884 12135 14886 12144
rect 14832 12106 14884 12112
rect 14844 11286 14872 12106
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14844 10062 14872 10678
rect 15120 10606 15148 11698
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11082 15332 11494
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15764 10674 15792 11290
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14922 8528 14978 8537
rect 14922 8463 14978 8472
rect 15028 8480 15056 10066
rect 15120 9994 15148 10542
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 10266 15424 10406
rect 15764 10266 15792 10610
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15396 10062 15424 10202
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 9178 15332 9454
rect 15764 9382 15792 10202
rect 15856 10062 15884 10542
rect 16408 10062 16436 12378
rect 16960 12238 16988 13806
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 11694 16988 12174
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16684 11354 16712 11630
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16776 11082 16804 11630
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 15856 9518 15884 9998
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9722 16436 9862
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9586 16528 10950
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 9654 16620 10406
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16684 9722 16712 9998
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15396 9178 15424 9318
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15396 8974 15424 9114
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15764 8838 15792 9046
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14476 7398 14780 7426
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13188 5302 13216 5646
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13556 4758 13584 6326
rect 13832 6066 13860 6734
rect 14384 6730 14412 7142
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 13740 6038 13860 6066
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13740 5914 13768 6038
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13740 5098 13768 5850
rect 13832 5234 13860 5850
rect 13924 5846 13952 6054
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 14108 5710 14136 6054
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14200 5642 14228 6666
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13544 4752 13596 4758
rect 13924 4729 13952 5170
rect 13544 4694 13596 4700
rect 13910 4720 13966 4729
rect 12992 4684 13044 4690
rect 13910 4655 13966 4664
rect 12992 4626 13044 4632
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12768 4168 12940 4196
rect 12716 4150 12768 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 3738 12664 4082
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12716 3664 12768 3670
rect 12452 3612 12716 3618
rect 12452 3606 12768 3612
rect 12452 3590 12756 3606
rect 12452 3516 12480 3590
rect 12360 3488 12480 3516
rect 12530 3496 12586 3505
rect 12164 3470 12216 3476
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11992 2854 12020 3402
rect 12176 3126 12204 3470
rect 12530 3431 12586 3440
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12084 2650 12112 2994
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 11428 1896 11480 1902
rect 11428 1838 11480 1844
rect 11796 1148 11848 1154
rect 11796 1090 11848 1096
rect 11808 800 11836 1090
rect 12176 800 12204 1974
rect 12544 800 12572 3431
rect 12912 2446 12940 3878
rect 13188 3058 13216 4558
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 13464 3534 13492 4422
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13188 2854 13216 2994
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13266 2544 13322 2553
rect 13266 2479 13322 2488
rect 12900 2440 12952 2446
rect 12806 2408 12862 2417
rect 12900 2382 12952 2388
rect 12806 2343 12862 2352
rect 12820 1170 12848 2343
rect 12820 1142 12940 1170
rect 12912 800 12940 1142
rect 13280 800 13308 2479
rect 13648 800 13676 3130
rect 13740 3058 13768 4218
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13910 3768 13966 3777
rect 13910 3703 13966 3712
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13832 2938 13860 3538
rect 13924 3126 13952 3703
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13832 2910 13952 2938
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2378 13860 2790
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13924 1850 13952 2910
rect 14016 2514 14044 3878
rect 14200 3194 14228 4082
rect 14292 4078 14320 4422
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 14108 2650 14136 2858
rect 14292 2854 14320 4014
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14372 2100 14424 2106
rect 14372 2042 14424 2048
rect 13924 1822 14044 1850
rect 14016 800 14044 1822
rect 14384 800 14412 2042
rect 10704 734 10916 762
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14476 762 14504 7398
rect 14844 6662 14872 8298
rect 14936 7410 14964 8463
rect 15028 8452 15148 8480
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14660 6322 14688 6598
rect 14936 6322 14964 7210
rect 15028 6798 15056 8298
rect 15120 8090 15148 8452
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15120 7546 15148 7686
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14568 5370 14596 6258
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14660 4826 14688 6258
rect 15120 5914 15148 6666
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14752 3738 14780 5714
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14752 3058 14780 3674
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14844 2446 14872 5646
rect 14936 5370 14964 5850
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15028 4622 15056 5578
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15120 4162 15148 5510
rect 15304 5409 15332 8774
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 7410 15424 8026
rect 15488 7750 15516 8434
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 8090 15608 8230
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15488 7342 15516 7686
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15580 6458 15608 7346
rect 15856 7206 15884 8910
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16316 8362 16344 8570
rect 16500 8498 16528 9522
rect 16776 8974 16804 11018
rect 16868 10266 16896 11562
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16960 10470 16988 10610
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16948 9580 17000 9586
rect 16868 9540 16948 9568
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 7410 15976 7822
rect 15936 7404 15988 7410
rect 15988 7364 16068 7392
rect 15936 7346 15988 7352
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 16040 6458 16068 7364
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6934 16252 7142
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15856 5710 15884 5850
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15290 5400 15346 5409
rect 15290 5335 15346 5344
rect 16040 5302 16068 6394
rect 16316 5846 16344 8298
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16408 6934 16436 7414
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16684 6882 16712 8366
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7478 16804 8230
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16684 6854 16804 6882
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6458 16712 6734
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16316 5574 16344 5782
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15028 4134 15148 4162
rect 14922 4040 14978 4049
rect 15028 4010 15056 4134
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14922 3975 14978 3984
rect 15016 4004 15068 4010
rect 14936 3126 14964 3975
rect 15016 3946 15068 3952
rect 15014 3224 15070 3233
rect 15014 3159 15070 3168
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15028 2530 15056 3159
rect 15120 2990 15148 4014
rect 15212 3534 15240 5238
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15474 4856 15530 4865
rect 15474 4791 15530 4800
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15304 4214 15332 4558
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15304 3058 15332 4150
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 14936 2502 15056 2530
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14936 1850 14964 2502
rect 15016 2440 15068 2446
rect 15120 2428 15148 2926
rect 15304 2446 15332 2994
rect 15068 2400 15148 2428
rect 15292 2440 15344 2446
rect 15016 2382 15068 2388
rect 15292 2382 15344 2388
rect 14936 1822 15148 1850
rect 14660 870 14780 898
rect 14660 762 14688 870
rect 14752 800 14780 870
rect 15120 800 15148 1822
rect 15488 800 15516 4791
rect 15948 4758 15976 5170
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 14476 734 14688 762
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15580 762 15608 4626
rect 16408 4622 16436 4966
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 4282 16436 4558
rect 16500 4554 16528 6054
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16776 4146 16804 6854
rect 16868 5137 16896 9540
rect 16948 9522 17000 9528
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 8498 16988 8570
rect 17144 8537 17172 13126
rect 17604 12714 17632 14282
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 19260 14006 19288 14214
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 20088 13938 20116 14418
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20272 13938 20300 14214
rect 20456 14074 20484 14350
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19444 13190 19472 13738
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12102 17448 12582
rect 17498 12200 17554 12209
rect 17498 12135 17500 12144
rect 17552 12135 17554 12144
rect 17500 12106 17552 12112
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17130 8528 17186 8537
rect 16948 8492 17000 8498
rect 17000 8452 17080 8480
rect 17130 8463 17186 8472
rect 16948 8434 17000 8440
rect 17052 7018 17080 8452
rect 17236 8294 17264 9454
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17052 6990 17172 7018
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16960 5846 16988 6258
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16854 5128 16910 5137
rect 16854 5063 16910 5072
rect 16960 4706 16988 5782
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 4826 17080 5170
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16960 4690 17080 4706
rect 16960 4684 17092 4690
rect 16960 4678 17040 4684
rect 17040 4626 17092 4632
rect 16120 4140 16172 4146
rect 16764 4140 16816 4146
rect 16120 4082 16172 4088
rect 16684 4100 16764 4128
rect 16132 3738 16160 4082
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16500 3534 16528 3878
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15764 2774 15792 3402
rect 16408 3058 16436 3470
rect 16684 3194 16712 4100
rect 16764 4082 16816 4088
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16776 3126 16804 3402
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 15764 2746 15884 2774
rect 15856 2650 15884 2746
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 16040 2446 16068 2790
rect 16776 2774 16804 3062
rect 16684 2746 16804 2774
rect 16684 2446 16712 2746
rect 16868 2446 16896 3878
rect 17052 2961 17080 4626
rect 17144 4622 17172 6990
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17236 3126 17264 6394
rect 17328 5846 17356 9522
rect 17420 7410 17448 10678
rect 17512 10538 17540 11698
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17604 10266 17632 12650
rect 17696 11014 17724 12786
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17972 11082 18000 12650
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 18248 12434 18276 12582
rect 19168 12442 19196 12582
rect 19156 12436 19208 12442
rect 18248 12406 18368 12434
rect 18050 12336 18106 12345
rect 18050 12271 18052 12280
rect 18104 12271 18106 12280
rect 18052 12242 18104 12248
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 11218 18184 11494
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10810 17724 10950
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 18064 10674 18092 11086
rect 18156 10742 18184 11154
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17604 8838 17632 10202
rect 17972 9994 18000 10202
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18064 9654 18092 9862
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17880 8974 17908 9454
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17880 8430 17908 8910
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17972 8090 18000 8434
rect 18064 8362 18092 8774
rect 18156 8362 18184 9998
rect 18248 9654 18276 11222
rect 18340 11150 18368 12406
rect 19156 12378 19208 12384
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18432 11218 18460 12310
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18432 10742 18460 11154
rect 18616 11150 18644 11562
rect 19168 11558 19196 12174
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18524 10538 18552 10746
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18340 9110 18368 10134
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17512 6118 17540 6938
rect 17880 6662 17908 7754
rect 17972 7546 18000 8026
rect 18064 7818 18092 8298
rect 18432 8090 18460 9862
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17972 6798 18000 7482
rect 18064 6866 18092 7754
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18248 6730 18276 7686
rect 18432 7002 18460 8026
rect 18524 7410 18552 10474
rect 18616 10266 18644 11086
rect 19168 10606 19196 11494
rect 19260 10810 19288 12854
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19168 10282 19196 10542
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18984 10254 19196 10282
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 7954 18644 8230
rect 18708 7954 18736 8298
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18800 7585 18828 10134
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18892 8090 18920 9114
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18328 6724 18380 6730
rect 18328 6666 18380 6672
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17604 5914 17632 6190
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17328 5710 17356 5782
rect 18248 5710 18276 6666
rect 18340 6186 18368 6666
rect 18432 6254 18460 6802
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18340 5642 18368 6122
rect 18432 5846 18460 6190
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18340 5370 18368 5578
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18340 4690 18368 5306
rect 18432 5302 18460 5782
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18432 4690 18460 5238
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17038 2952 17094 2961
rect 17038 2887 17094 2896
rect 17328 2582 17356 3402
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17316 2576 17368 2582
rect 17316 2518 17368 2524
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 15764 870 15884 898
rect 15764 762 15792 870
rect 15856 800 15884 870
rect 16592 800 16620 2314
rect 17420 800 17448 2518
rect 17788 2514 17816 3334
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17972 2446 18000 3946
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18156 800 18184 2790
rect 18248 2446 18276 3878
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18616 2106 18644 5510
rect 18708 2650 18736 6734
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18800 4826 18828 5170
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18892 4146 18920 7210
rect 18984 5710 19012 10254
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19168 8378 19196 8910
rect 19352 8566 19380 13126
rect 19444 12850 19472 13126
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19996 12850 20024 13194
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19996 12442 20024 12786
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20088 12170 20116 13262
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11150 19472 12038
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 9382 19472 11086
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19904 10470 19932 10542
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19996 9568 20024 11154
rect 19628 9540 20024 9568
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9081 19472 9318
rect 19430 9072 19486 9081
rect 19628 9042 19656 9540
rect 19996 9450 20024 9540
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19720 9353 19748 9386
rect 19706 9344 19762 9353
rect 19706 9279 19762 9288
rect 20180 9178 20208 13330
rect 20272 12782 20300 13874
rect 20732 13394 20760 14758
rect 21376 14414 21404 14758
rect 21928 14498 21956 14894
rect 22020 14618 22048 14962
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21928 14470 22048 14498
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21192 13870 21220 14350
rect 21376 14006 21404 14350
rect 22020 14278 22048 14470
rect 22204 14414 22232 14758
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21548 14000 21600 14006
rect 21836 13988 21864 14214
rect 21916 14000 21968 14006
rect 21836 13960 21916 13988
rect 21548 13942 21600 13948
rect 21916 13942 21968 13948
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20732 12238 20760 13330
rect 20824 12730 20852 13398
rect 20916 13326 20944 13398
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 12986 21036 13126
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20824 12702 21036 12730
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12232 20772 12238
rect 20534 12200 20590 12209
rect 20720 12174 20772 12180
rect 20534 12135 20536 12144
rect 20588 12135 20590 12144
rect 20536 12106 20588 12112
rect 20732 11830 20760 12174
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20548 11354 20576 11698
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20824 11150 20852 12582
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20350 10568 20406 10577
rect 20350 10503 20352 10512
rect 20404 10503 20406 10512
rect 20352 10474 20404 10480
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 9586 20484 10406
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20732 9586 20760 9658
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 19430 9007 19486 9016
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19904 9030 20116 9058
rect 19904 8906 19932 9030
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19168 8350 19380 8378
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7546 19104 7822
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6458 19288 6598
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19352 5846 19380 8350
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19064 5228 19116 5234
rect 19352 5216 19380 5782
rect 19064 5170 19116 5176
rect 19168 5188 19380 5216
rect 19076 4622 19104 5170
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 4214 19104 4558
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 19076 3126 19104 4150
rect 19168 4146 19196 5188
rect 19444 5114 19472 8774
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19904 7993 19932 8502
rect 19996 8498 20024 8910
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19890 7984 19946 7993
rect 19890 7919 19946 7928
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19536 6644 19564 7414
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 19720 6798 19748 6870
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19516 6616 19564 6644
rect 19516 6440 19544 6616
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19996 6458 20024 7346
rect 19984 6452 20036 6458
rect 19516 6412 19564 6440
rect 19536 5710 19564 6412
rect 19984 6394 20036 6400
rect 20088 6338 20116 9030
rect 20364 8974 20392 9279
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20180 8634 20208 8910
rect 20456 8906 20484 9522
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20166 8120 20222 8129
rect 20166 8055 20222 8064
rect 20180 7478 20208 8055
rect 20168 7472 20220 7478
rect 20168 7414 20220 7420
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19996 6310 20116 6338
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19352 5086 19472 5114
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19168 3058 19196 3878
rect 19260 3602 19288 4626
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19352 3534 19380 5086
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 19444 2446 19472 4966
rect 19996 4622 20024 6310
rect 20180 5710 20208 7278
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6390 20300 7142
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20272 5234 20300 6122
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 2446 20024 4422
rect 20088 4146 20116 5034
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 4282 20208 4422
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20364 2990 20392 8774
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20456 4554 20484 8434
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7206 20576 7686
rect 20640 7478 20668 9386
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 5914 20576 7142
rect 20640 6254 20668 7414
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20548 5370 20576 5714
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20640 4826 20668 5578
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20456 3194 20484 4490
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20640 3058 20668 3334
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20732 2446 20760 4966
rect 20824 4622 20852 9114
rect 20916 6730 20944 11018
rect 21008 9704 21036 12702
rect 21100 12170 21128 13670
rect 21192 12434 21220 13806
rect 21192 12406 21312 12434
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21192 11898 21220 12106
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21192 10266 21220 10610
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21008 9676 21220 9704
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 9110 21036 9522
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21100 9042 21128 9386
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20996 7880 21048 7886
rect 21192 7868 21220 9676
rect 21284 8974 21312 12406
rect 21376 12238 21404 13942
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11558 21404 12038
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 10742 21404 11494
rect 21468 10742 21496 13806
rect 21560 13462 21588 13942
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21560 12102 21588 13398
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21652 12850 21680 13330
rect 21732 13320 21784 13326
rect 21928 13308 21956 13942
rect 22020 13870 22048 14214
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 21784 13280 21956 13308
rect 21732 13262 21784 13268
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21744 12238 21772 12378
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21376 8498 21404 10678
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21272 7880 21324 7886
rect 21192 7840 21272 7868
rect 20996 7822 21048 7828
rect 21272 7822 21324 7828
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20902 5672 20958 5681
rect 20902 5607 20904 5616
rect 20956 5607 20958 5616
rect 20904 5578 20956 5584
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20916 3194 20944 5102
rect 21008 4554 21036 7822
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21192 7002 21220 7686
rect 21284 7410 21312 7686
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21468 6186 21496 7210
rect 21560 6390 21588 7754
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21008 4214 21036 4490
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 21100 4146 21128 4558
rect 21652 4146 21680 12174
rect 21744 8786 21772 12174
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11626 21864 12038
rect 21928 11694 21956 13280
rect 22020 13190 22048 13670
rect 22296 13530 22324 13670
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22020 11898 22048 13126
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22112 11762 22140 13126
rect 22296 12782 22324 13466
rect 22388 12986 22416 13874
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22664 12646 22692 15642
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22848 15162 22876 15302
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 23032 14414 23060 15030
rect 23400 14618 23428 15370
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23032 13870 23060 14350
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22756 12170 22784 13806
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22388 11898 22416 12106
rect 22940 11898 22968 13194
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21836 9722 21864 10610
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21744 8758 21864 8786
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21744 7818 21772 8570
rect 21836 7954 21864 8758
rect 21928 8498 21956 9318
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21560 3738 21588 4014
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21744 3534 21772 7754
rect 21824 7540 21876 7546
rect 21928 7528 21956 7754
rect 21876 7500 21956 7528
rect 21824 7482 21876 7488
rect 22020 7342 22048 11562
rect 22112 10674 22140 11698
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22100 9648 22152 9654
rect 22098 9616 22100 9625
rect 22152 9616 22154 9625
rect 22098 9551 22154 9560
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 21928 7154 21956 7210
rect 22204 7154 22232 11086
rect 22296 9586 22324 11766
rect 23032 11762 23060 13806
rect 23308 12306 23336 14486
rect 23492 13802 23520 15914
rect 23584 15348 23612 16186
rect 23676 15502 23704 16390
rect 23768 15502 23796 16526
rect 25148 16182 25176 16526
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23664 15360 23716 15366
rect 23584 15320 23664 15348
rect 23664 15302 23716 15308
rect 23676 13870 23704 15302
rect 23860 15026 23888 15846
rect 24320 15706 24348 16050
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 25148 15502 25176 16118
rect 26252 16114 26280 16390
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26252 15994 26280 16050
rect 26700 16040 26752 16046
rect 26252 15966 26372 15994
rect 26700 15982 26752 15988
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 24964 15162 24992 15438
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22296 9042 22324 9522
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 8650 22324 8842
rect 22388 8838 22416 11154
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 9586 22508 10474
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22572 8906 22600 11494
rect 23676 11354 23704 11698
rect 23768 11694 23796 13126
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22296 8622 22600 8650
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22376 8492 22428 8498
rect 21928 7126 22232 7154
rect 22296 8452 22376 8480
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21928 5914 21956 6734
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 22296 5234 22324 8452
rect 22376 8434 22428 8440
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21008 3058 21036 3402
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21836 2990 21864 4422
rect 22112 4146 22140 5170
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22204 4146 22232 5102
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22204 3466 22232 3946
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18892 800 18920 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 898 20024 2246
rect 19628 870 19748 898
rect 19628 800 19656 870
rect 15580 734 15792 762
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19720 762 19748 870
rect 19904 870 20024 898
rect 19904 762 19932 870
rect 20364 800 20392 2246
rect 21100 800 21128 2518
rect 21836 800 21864 2790
rect 22204 2650 22232 3402
rect 22388 3058 22416 8298
rect 22480 7546 22508 8502
rect 22572 8242 22600 8622
rect 22664 8362 22692 9930
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22756 9489 22784 9590
rect 22742 9480 22798 9489
rect 22742 9415 22798 9424
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22756 8242 22784 8842
rect 22848 8566 22876 10746
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 22572 8214 22784 8242
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22480 7410 22508 7482
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22572 6934 22600 8214
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 7002 22692 7346
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22560 6928 22612 6934
rect 22560 6870 22612 6876
rect 22652 6792 22704 6798
rect 22572 6752 22652 6780
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22480 6458 22508 6598
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22480 5522 22508 6394
rect 22572 6322 22600 6752
rect 22652 6734 22704 6740
rect 22756 6662 22784 7278
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22572 5817 22600 6258
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22558 5808 22614 5817
rect 22558 5743 22560 5752
rect 22612 5743 22614 5752
rect 22560 5714 22612 5720
rect 22480 5494 22600 5522
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22480 4690 22508 5306
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22480 3738 22508 4626
rect 22572 4622 22600 5494
rect 22664 5302 22692 6054
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22572 800 22600 3878
rect 22664 2378 22692 4218
rect 22848 3534 22876 8298
rect 22940 7002 22968 10406
rect 23032 10062 23060 11086
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22926 6488 22982 6497
rect 22926 6423 22982 6432
rect 22940 6390 22968 6423
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23032 5778 23060 9998
rect 23124 8430 23152 10610
rect 23216 10470 23244 11018
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23032 5370 23060 5714
rect 23124 5574 23152 6666
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 22928 5092 22980 5098
rect 22928 5034 22980 5040
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22940 2446 22968 5034
rect 23032 4622 23060 5306
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23124 2854 23152 5306
rect 23216 5114 23244 10406
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7410 23428 7686
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23400 7274 23428 7346
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23308 5234 23336 7142
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23216 5086 23336 5114
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23216 3602 23244 4014
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23216 3058 23244 3538
rect 23308 3058 23336 5086
rect 23400 4706 23428 6054
rect 23492 5234 23520 10406
rect 23584 9178 23612 10678
rect 23860 10674 23888 14962
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24308 14408 24360 14414
rect 24412 14362 24440 14758
rect 24780 14618 24808 14758
rect 25424 14618 25452 15030
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25608 14414 25636 15302
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 25872 14544 25924 14550
rect 25872 14486 25924 14492
rect 25884 14414 25912 14486
rect 24360 14356 24440 14362
rect 24308 14350 24440 14356
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 24320 14334 24440 14350
rect 24412 13938 24440 14334
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24228 12986 24256 13874
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24412 12306 24440 13874
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 12374 24532 13806
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24492 12368 24544 12374
rect 24492 12310 24544 12316
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24308 11280 24360 11286
rect 24308 11222 24360 11228
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23952 10577 23980 10678
rect 23938 10568 23994 10577
rect 23938 10503 23994 10512
rect 24216 10532 24268 10538
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23768 9722 23796 9930
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23754 9616 23810 9625
rect 23754 9551 23810 9560
rect 23768 9518 23796 9551
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23570 9072 23626 9081
rect 23570 9007 23626 9016
rect 23584 8498 23612 9007
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23676 7970 23704 8502
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23584 7942 23704 7970
rect 23584 7274 23612 7942
rect 23768 7886 23796 8434
rect 23860 8090 23888 8434
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23584 7002 23612 7210
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23676 6254 23704 7822
rect 23952 7410 23980 10503
rect 24216 10474 24268 10480
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 9042 24072 9522
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 23952 6866 23980 7346
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 6180 23624 6186
rect 23572 6122 23624 6128
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23400 4678 23520 4706
rect 23386 4584 23442 4593
rect 23386 4519 23388 4528
rect 23440 4519 23442 4528
rect 23388 4490 23440 4496
rect 23492 4434 23520 4678
rect 23400 4406 23520 4434
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 23400 800 23428 4406
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3738 23520 4082
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23584 3194 23612 6122
rect 23676 5710 23704 6190
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 24136 5234 24164 7686
rect 24228 6322 24256 10474
rect 24320 9654 24348 11222
rect 24504 9874 24532 12310
rect 24596 12170 24624 12922
rect 24780 12442 24808 14214
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24872 13326 24900 13806
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24964 12442 24992 13330
rect 25056 13258 25084 14350
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 13938 25176 14282
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24596 10062 24624 12106
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24688 11354 24716 11698
rect 25056 11354 25084 13194
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25148 11150 25176 13874
rect 25332 12850 25360 14214
rect 25608 14006 25636 14350
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25608 11830 25636 12174
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25976 12050 26004 13942
rect 26068 12170 26096 14758
rect 26160 13734 26188 14826
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26344 13954 26372 15966
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26436 14074 26464 14962
rect 26712 14958 26740 15982
rect 26988 15978 27016 16458
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 26976 15972 27028 15978
rect 26976 15914 27028 15920
rect 27172 15502 27200 16390
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27816 15162 27844 16526
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28368 16114 28396 16390
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28828 15638 28856 16526
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28920 15706 28948 16458
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29104 15892 29132 16390
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 29184 15904 29236 15910
rect 29104 15864 29184 15892
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 28816 15632 28868 15638
rect 28816 15574 28868 15580
rect 27896 15360 27948 15366
rect 27896 15302 27948 15308
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27344 15088 27396 15094
rect 27344 15030 27396 15036
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26712 14618 26740 14894
rect 27356 14618 27384 15030
rect 27908 15026 27936 15302
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26160 12850 26188 13330
rect 26252 12986 26280 13942
rect 26344 13926 26464 13954
rect 26436 13190 26464 13926
rect 26528 13870 26556 14350
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26528 13326 26556 13806
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26344 12782 26372 13126
rect 26436 12850 26464 13126
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26528 12714 26556 13262
rect 27344 13184 27396 13190
rect 27344 13126 27396 13132
rect 27356 12850 27384 13126
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 26884 12776 26936 12782
rect 26884 12718 26936 12724
rect 26516 12708 26568 12714
rect 26516 12650 26568 12656
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 26896 12084 26924 12718
rect 26988 12434 27016 12786
rect 26988 12406 27292 12434
rect 27160 12368 27212 12374
rect 27160 12310 27212 12316
rect 26976 12096 27028 12102
rect 26896 12056 26976 12084
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25136 11144 25188 11150
rect 25188 11092 25360 11098
rect 25136 11086 25360 11092
rect 25148 11082 25360 11086
rect 25700 11082 25728 12038
rect 25976 12022 26096 12050
rect 26976 12038 27028 12044
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25148 11076 25372 11082
rect 25148 11070 25320 11076
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24504 9846 24624 9874
rect 24308 9648 24360 9654
rect 24308 9590 24360 9596
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24412 6866 24440 7414
rect 24596 6866 24624 9846
rect 24688 9722 24716 10610
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24676 9716 24728 9722
rect 24872 9704 24900 9998
rect 25056 9926 25084 10950
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 24676 9658 24728 9664
rect 24780 9676 24900 9704
rect 24688 8498 24716 9658
rect 24780 9178 24808 9676
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24780 8566 24808 9114
rect 24872 9110 24900 9522
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24964 8498 24992 9862
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24688 7818 24716 8434
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24766 8120 24822 8129
rect 24766 8055 24768 8064
rect 24820 8055 24822 8064
rect 24768 8026 24820 8032
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24688 6798 24716 7754
rect 24872 7546 24900 8298
rect 25056 8106 25084 9862
rect 24964 8078 25084 8106
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24872 6798 24900 7346
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23860 4826 23888 5170
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23952 4622 23980 5034
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23952 4146 23980 4558
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 24412 3942 24440 5034
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 24596 3058 24624 6598
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24872 4146 24900 4490
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24964 3534 24992 8078
rect 25148 7342 25176 11070
rect 25320 11018 25372 11024
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25792 11014 25820 11494
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25884 11150 25912 11290
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25240 8838 25268 9454
rect 25332 8838 25360 9998
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25424 9722 25452 9930
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25318 7984 25374 7993
rect 25318 7919 25320 7928
rect 25372 7919 25374 7928
rect 25320 7890 25372 7896
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25148 6254 25176 6734
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25228 6180 25280 6186
rect 25228 6122 25280 6128
rect 25240 4570 25268 6122
rect 25424 5681 25452 9318
rect 25516 8673 25544 10406
rect 25608 10130 25636 10610
rect 25688 10464 25740 10470
rect 25884 10418 25912 10950
rect 25688 10406 25740 10412
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25608 9722 25636 10066
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 25502 8664 25558 8673
rect 25502 8599 25558 8608
rect 25594 8528 25650 8537
rect 25594 8463 25596 8472
rect 25648 8463 25650 8472
rect 25596 8434 25648 8440
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25516 7886 25544 8298
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25410 5672 25466 5681
rect 25410 5607 25466 5616
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4622 25452 4966
rect 25056 4542 25268 4570
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24872 3058 24900 3334
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 24136 800 24164 2246
rect 24872 800 24900 2790
rect 25056 2446 25084 4542
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25148 4078 25176 4422
rect 25424 4282 25452 4558
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25148 2446 25176 4014
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 25240 2854 25268 3402
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25516 2514 25544 7822
rect 25608 7410 25636 8230
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25608 7206 25636 7346
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25608 6798 25636 7142
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25700 5642 25728 10406
rect 25792 10390 25912 10418
rect 25792 8090 25820 10390
rect 26068 10180 26096 12022
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 25976 10152 26096 10180
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25884 9586 25912 9998
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25976 8922 26004 10152
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 26068 9586 26096 9862
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26160 9042 26188 11154
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 25976 8894 26188 8922
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25688 5636 25740 5642
rect 25688 5578 25740 5584
rect 25780 4208 25832 4214
rect 25780 4150 25832 4156
rect 25792 4078 25820 4150
rect 25884 4128 25912 8774
rect 25976 8566 26004 8774
rect 25964 8560 26016 8566
rect 25964 8502 26016 8508
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25976 5846 26004 6054
rect 26068 5914 26096 7278
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 25964 5840 26016 5846
rect 25964 5782 26016 5788
rect 26056 4548 26108 4554
rect 26056 4490 26108 4496
rect 26068 4282 26096 4490
rect 26056 4276 26108 4282
rect 26056 4218 26108 4224
rect 25962 4176 26018 4185
rect 26160 4146 26188 8894
rect 26252 5642 26280 11494
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26344 8090 26372 9114
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 25884 4120 25962 4128
rect 25884 4100 25964 4120
rect 26016 4111 26018 4120
rect 26148 4140 26200 4146
rect 25964 4082 26016 4088
rect 26148 4082 26200 4088
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25792 3194 25820 4014
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25976 3058 26004 4082
rect 26344 3738 26372 6734
rect 26436 5370 26464 11698
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26528 7002 26556 10610
rect 26620 10470 26648 11766
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26896 11286 26924 11562
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 10130 26648 10406
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26620 9518 26648 10066
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26804 9042 26832 9590
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26606 8664 26662 8673
rect 26606 8599 26662 8608
rect 26620 8498 26648 8599
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26620 8090 26648 8434
rect 26712 8430 26740 8910
rect 26804 8430 26832 8978
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 26608 8084 26660 8090
rect 26608 8026 26660 8032
rect 26804 7478 26832 8366
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 26528 6390 26556 6938
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 26804 6254 26832 7210
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26528 5574 26556 6190
rect 26700 6180 26752 6186
rect 26700 6122 26752 6128
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 26436 4826 26464 5102
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 26528 2990 26556 5510
rect 26712 4826 26740 6122
rect 26896 5642 26924 6734
rect 26988 6322 27016 12038
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27080 11354 27108 11698
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27172 11150 27200 12310
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27080 6798 27108 7278
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27172 6458 27200 9522
rect 27264 8634 27292 12406
rect 27540 11830 27568 13262
rect 27632 12986 27660 13942
rect 27724 13938 27752 14350
rect 27816 14278 27844 14894
rect 27908 14346 27936 14962
rect 28828 14958 28856 15574
rect 29012 15570 29040 15846
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 29104 15502 29132 15864
rect 29184 15846 29236 15852
rect 30300 15706 30328 16050
rect 30760 15706 30788 16050
rect 31300 15904 31352 15910
rect 31300 15846 31352 15852
rect 31576 15904 31628 15910
rect 31576 15846 31628 15852
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 30748 15700 30800 15706
rect 30748 15642 30800 15648
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 28816 14952 28868 14958
rect 28736 14900 28816 14906
rect 28736 14894 28868 14900
rect 28736 14878 28856 14894
rect 28632 14816 28684 14822
rect 28632 14758 28684 14764
rect 28644 14414 28672 14758
rect 28736 14618 28764 14878
rect 28724 14612 28776 14618
rect 28724 14554 28776 14560
rect 28632 14408 28684 14414
rect 28632 14350 28684 14356
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27804 14272 27856 14278
rect 27804 14214 27856 14220
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27724 11354 27752 12174
rect 27816 12102 27844 14214
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27356 11014 27384 11086
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27908 10418 27936 14282
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 28000 14074 28028 14214
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 28356 14000 28408 14006
rect 28356 13942 28408 13948
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 28000 12782 28028 13874
rect 28368 12782 28396 13942
rect 28644 13938 28672 14350
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28920 14074 28948 14214
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28460 13190 28488 13874
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28644 12850 28672 13874
rect 29012 13326 29040 14214
rect 29104 14006 29132 15438
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30484 14618 30512 15370
rect 30668 15162 30696 15438
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 31128 14482 31156 15506
rect 31312 15502 31340 15846
rect 31300 15496 31352 15502
rect 31300 15438 31352 15444
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30380 14408 30432 14414
rect 30380 14350 30432 14356
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28000 12238 28028 12718
rect 28736 12714 28764 13126
rect 29000 12844 29052 12850
rect 29104 12832 29132 13942
rect 29656 13938 29684 14214
rect 29748 14074 29776 14350
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29288 13462 29316 13806
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29276 13456 29328 13462
rect 29276 13398 29328 13404
rect 29564 13394 29592 13670
rect 29552 13388 29604 13394
rect 29552 13330 29604 13336
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29840 12850 29868 13330
rect 29052 12804 29132 12832
rect 29828 12844 29880 12850
rect 29000 12786 29052 12792
rect 29828 12786 29880 12792
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 28724 12708 28776 12714
rect 28724 12650 28776 12656
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 27724 10390 27936 10418
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27540 8537 27568 8910
rect 27526 8528 27582 8537
rect 27724 8498 27752 10390
rect 27526 8463 27528 8472
rect 27580 8463 27582 8472
rect 27712 8492 27764 8498
rect 27528 8434 27580 8440
rect 27712 8434 27764 8440
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27356 6866 27384 7482
rect 27448 7478 27476 7822
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27448 7002 27476 7414
rect 27540 7002 27568 7686
rect 27908 7546 27936 8434
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28000 7426 28028 8298
rect 27908 7398 28028 7426
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27356 6322 27384 6802
rect 27908 6798 27936 7398
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 27986 6760 28042 6769
rect 27448 6390 27476 6734
rect 27620 6724 27672 6730
rect 27620 6666 27672 6672
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 26976 6316 27028 6322
rect 26976 6258 27028 6264
rect 27344 6316 27396 6322
rect 27344 6258 27396 6264
rect 27448 6202 27476 6326
rect 27264 6174 27476 6202
rect 27264 5710 27292 6174
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27342 5944 27398 5953
rect 27342 5879 27398 5888
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 26884 5636 26936 5642
rect 26884 5578 26936 5584
rect 26896 5166 26924 5578
rect 27264 5234 27292 5646
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26804 4826 26832 4966
rect 26700 4820 26752 4826
rect 26700 4762 26752 4768
rect 26792 4820 26844 4826
rect 26792 4762 26844 4768
rect 27356 4146 27384 5879
rect 27448 5370 27476 6054
rect 27632 5846 27660 6666
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27816 5914 27844 6394
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27632 5386 27660 5782
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27540 5358 27660 5386
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 26804 3738 26832 4082
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 27342 3496 27398 3505
rect 27342 3431 27344 3440
rect 27396 3431 27398 3440
rect 27344 3402 27396 3408
rect 27448 3058 27476 5306
rect 27540 5030 27568 5358
rect 27620 5296 27672 5302
rect 27620 5238 27672 5244
rect 27712 5296 27764 5302
rect 27712 5238 27764 5244
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27540 4622 27568 4966
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27540 4486 27568 4558
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27540 4282 27568 4422
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 27528 3528 27580 3534
rect 27632 3516 27660 5238
rect 27724 4690 27752 5238
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27816 4146 27844 5510
rect 27804 4140 27856 4146
rect 27580 3488 27660 3516
rect 27724 4100 27804 4128
rect 27528 3470 27580 3476
rect 27724 3058 27752 4100
rect 27804 4082 27856 4088
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 27068 2916 27120 2922
rect 27068 2858 27120 2864
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25608 800 25636 2518
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26344 800 26372 2246
rect 27080 800 27108 2858
rect 27816 800 27844 3130
rect 27908 3058 27936 6734
rect 27986 6695 27988 6704
rect 28040 6695 28042 6704
rect 27988 6666 28040 6672
rect 28092 6322 28120 12650
rect 29012 12646 29040 12786
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29656 12434 29684 12582
rect 29656 12406 29776 12434
rect 28630 12200 28686 12209
rect 28630 12135 28632 12144
rect 28684 12135 28686 12144
rect 28632 12106 28684 12112
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28276 11558 28304 12038
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28276 11218 28304 11494
rect 28644 11354 28672 12106
rect 29644 12096 29696 12102
rect 29644 12038 29696 12044
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28184 8634 28212 9046
rect 28276 8974 28304 11154
rect 28908 11144 28960 11150
rect 29012 11098 29040 11834
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 28960 11092 29040 11098
rect 28908 11086 29040 11092
rect 28920 11070 29040 11086
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28368 10044 28396 10746
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 28460 10198 28488 10678
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 28920 10266 28948 10610
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28448 10192 28500 10198
rect 28448 10134 28500 10140
rect 28448 10056 28500 10062
rect 28368 10016 28448 10044
rect 28448 9998 28500 10004
rect 28632 10056 28684 10062
rect 28632 9998 28684 10004
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 8974 28488 9862
rect 28264 8968 28316 8974
rect 28264 8910 28316 8916
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28184 8498 28212 8570
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28446 8256 28502 8265
rect 28446 8191 28502 8200
rect 28460 8090 28488 8191
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28184 6202 28212 7958
rect 28276 7868 28304 8026
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28356 7880 28408 7886
rect 28276 7840 28356 7868
rect 28356 7822 28408 7828
rect 28460 7818 28488 7890
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28552 7750 28580 8026
rect 28540 7744 28592 7750
rect 28540 7686 28592 7692
rect 28644 7206 28672 9998
rect 29012 9500 29040 11070
rect 29564 10674 29592 11494
rect 29656 10674 29684 12038
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 29104 9654 29132 10474
rect 29656 9994 29684 10610
rect 29644 9988 29696 9994
rect 29644 9930 29696 9936
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29092 9648 29144 9654
rect 29092 9590 29144 9596
rect 28722 9480 28778 9489
rect 29012 9472 29132 9500
rect 28722 9415 28724 9424
rect 28776 9415 28778 9424
rect 28724 9386 28776 9392
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 28724 9104 28776 9110
rect 28724 9046 28776 9052
rect 28736 8022 28764 9046
rect 28828 8498 28856 9114
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 28920 8498 28948 8842
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 28954 8356 29006 8362
rect 28954 8298 29006 8304
rect 28814 8256 28870 8265
rect 28966 8242 28994 8298
rect 28870 8214 28994 8242
rect 28814 8191 28870 8200
rect 28814 8120 28870 8129
rect 28814 8055 28870 8064
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28828 7954 28856 8055
rect 28998 7984 29054 7993
rect 28816 7948 28868 7954
rect 28998 7919 29054 7928
rect 28816 7890 28868 7896
rect 29012 7546 29040 7919
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28540 6792 28592 6798
rect 28540 6734 28592 6740
rect 28264 6724 28316 6730
rect 28264 6666 28316 6672
rect 28276 6497 28304 6666
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 28262 6488 28318 6497
rect 28262 6423 28318 6432
rect 28264 6316 28316 6322
rect 28264 6258 28316 6264
rect 28000 6174 28212 6202
rect 28000 4146 28028 6174
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28092 4826 28120 5646
rect 28170 5536 28226 5545
rect 28170 5471 28226 5480
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 27988 3460 28040 3466
rect 27988 3402 28040 3408
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 28000 2990 28028 3402
rect 27988 2984 28040 2990
rect 27988 2926 28040 2932
rect 28092 2650 28120 4626
rect 28184 3720 28212 5471
rect 28276 5370 28304 6258
rect 28460 6186 28488 6598
rect 28552 6322 28580 6734
rect 28540 6316 28592 6322
rect 28540 6258 28592 6264
rect 28448 6180 28500 6186
rect 28448 6122 28500 6128
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28368 4622 28396 6054
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28552 5098 28580 5646
rect 28540 5092 28592 5098
rect 28540 5034 28592 5040
rect 28644 4622 28672 7142
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 29012 5642 29040 6394
rect 29000 5636 29052 5642
rect 29000 5578 29052 5584
rect 29012 4622 29040 5578
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 28264 4548 28316 4554
rect 28264 4490 28316 4496
rect 28276 4146 28304 4490
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28264 3732 28316 3738
rect 28184 3692 28264 3720
rect 28264 3674 28316 3680
rect 28172 3528 28224 3534
rect 28170 3496 28172 3505
rect 28224 3496 28226 3505
rect 28170 3431 28226 3440
rect 28172 3120 28224 3126
rect 28224 3068 28304 3074
rect 28172 3062 28304 3068
rect 28184 3046 28304 3062
rect 28368 3058 28396 4558
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28170 2952 28226 2961
rect 28276 2938 28304 3046
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28276 2910 28396 2938
rect 28170 2887 28226 2896
rect 28184 2854 28212 2887
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28368 2650 28396 2910
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 28460 2514 28488 4422
rect 28724 4276 28776 4282
rect 28724 4218 28776 4224
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28540 2848 28592 2854
rect 28540 2790 28592 2796
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 28552 800 28580 2790
rect 28644 2378 28672 3878
rect 28736 3602 28764 4218
rect 28816 4208 28868 4214
rect 28816 4150 28868 4156
rect 28906 4176 28962 4185
rect 28828 3670 28856 4150
rect 28906 4111 28908 4120
rect 28960 4111 28962 4120
rect 28908 4082 28960 4088
rect 29012 4010 29040 4218
rect 29104 4146 29132 9472
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29196 8566 29224 9318
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29276 8356 29328 8362
rect 29276 8298 29328 8304
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29288 7818 29316 8298
rect 29276 7812 29328 7818
rect 29276 7754 29328 7760
rect 29288 6202 29316 7754
rect 29380 6322 29408 8298
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29288 6174 29408 6202
rect 29276 5228 29328 5234
rect 29196 5188 29276 5216
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 28724 3596 28776 3602
rect 28724 3538 28776 3544
rect 28828 2990 28856 3606
rect 29196 3466 29224 5188
rect 29276 5170 29328 5176
rect 29380 4729 29408 6174
rect 29472 4826 29500 9658
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29656 9042 29684 9318
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 29656 6390 29684 8978
rect 29748 6798 29776 12406
rect 29840 11150 29868 12786
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29932 12238 29960 12582
rect 30208 12442 30236 14350
rect 30392 13870 30420 14350
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30932 13864 30984 13870
rect 30932 13806 30984 13812
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30760 13462 30788 13670
rect 30748 13456 30800 13462
rect 30748 13398 30800 13404
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12646 30328 13194
rect 30760 13002 30788 13398
rect 30668 12974 30788 13002
rect 30944 12986 30972 13806
rect 31128 13802 31156 14418
rect 31312 14006 31340 15438
rect 31588 15094 31616 15846
rect 31944 15700 31996 15706
rect 31944 15642 31996 15648
rect 31576 15088 31628 15094
rect 31576 15030 31628 15036
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31404 14346 31432 14962
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31392 14340 31444 14346
rect 31392 14282 31444 14288
rect 31300 14000 31352 14006
rect 31300 13942 31352 13948
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 31116 13796 31168 13802
rect 31116 13738 31168 13744
rect 30932 12980 30984 12986
rect 30668 12918 30696 12974
rect 30932 12922 30984 12928
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 31024 12912 31076 12918
rect 31024 12854 31076 12860
rect 30288 12640 30340 12646
rect 30288 12582 30340 12588
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 29932 11218 29960 12174
rect 30668 12170 30696 12854
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30576 11830 30604 12038
rect 30564 11824 30616 11830
rect 30564 11766 30616 11772
rect 30760 11354 30788 12174
rect 31036 11898 31064 12854
rect 31128 12306 31156 13738
rect 31220 13326 31248 13874
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31404 13190 31432 14282
rect 31496 14074 31524 14350
rect 31588 14278 31616 15030
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31760 14272 31812 14278
rect 31760 14214 31812 14220
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31208 13184 31260 13190
rect 31208 13126 31260 13132
rect 31392 13184 31444 13190
rect 31392 13126 31444 13132
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31220 12918 31248 13126
rect 31404 12986 31432 13126
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 31208 12912 31260 12918
rect 31208 12854 31260 12860
rect 31496 12850 31524 13126
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31484 12844 31536 12850
rect 31484 12786 31536 12792
rect 31116 12300 31168 12306
rect 31116 12242 31168 12248
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31024 11892 31076 11898
rect 31024 11834 31076 11840
rect 30932 11688 30984 11694
rect 30932 11630 30984 11636
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 29840 10062 29868 11086
rect 30564 11008 30616 11014
rect 30564 10950 30616 10956
rect 30576 10742 30604 10950
rect 30564 10736 30616 10742
rect 30564 10678 30616 10684
rect 30564 10532 30616 10538
rect 30564 10474 30616 10480
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 30378 9888 30434 9897
rect 30378 9823 30434 9832
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 30024 8294 30052 8570
rect 30392 8294 30420 9823
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30484 8498 30512 8774
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30576 8430 30604 10474
rect 30668 10266 30696 11086
rect 30944 11014 30972 11630
rect 31220 11626 31248 12174
rect 31208 11620 31260 11626
rect 31208 11562 31260 11568
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30944 10810 30972 10950
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30760 10062 30788 10406
rect 30852 10130 30880 10406
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30012 8288 30064 8294
rect 30012 8230 30064 8236
rect 30380 8288 30432 8294
rect 30668 8242 30696 9862
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30760 8430 30788 8842
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 30380 8230 30432 8236
rect 30024 8022 30052 8230
rect 30012 8016 30064 8022
rect 30012 7958 30064 7964
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29644 6384 29696 6390
rect 29644 6326 29696 6332
rect 29840 5778 29868 7346
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 30208 6458 30236 6734
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 29828 5772 29880 5778
rect 29828 5714 29880 5720
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29644 4820 29696 4826
rect 29644 4762 29696 4768
rect 29366 4720 29422 4729
rect 29366 4655 29422 4664
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 29288 3738 29316 4082
rect 29276 3732 29328 3738
rect 29276 3674 29328 3680
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 29276 3596 29328 3602
rect 29380 3584 29408 3674
rect 29328 3556 29408 3584
rect 29276 3538 29328 3544
rect 29184 3460 29236 3466
rect 29184 3402 29236 3408
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 29000 2916 29052 2922
rect 29000 2858 29052 2864
rect 29012 2650 29040 2858
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29288 2582 29316 2790
rect 29276 2576 29328 2582
rect 29276 2518 29328 2524
rect 29368 2576 29420 2582
rect 29368 2518 29420 2524
rect 28632 2372 28684 2378
rect 28632 2314 28684 2320
rect 29380 800 29408 2518
rect 29564 2446 29592 4422
rect 29656 4214 29684 4762
rect 29828 4684 29880 4690
rect 29828 4626 29880 4632
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 29644 4208 29696 4214
rect 29644 4150 29696 4156
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 29656 2514 29684 3878
rect 29748 3058 29776 4422
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 29840 2990 29868 4626
rect 29828 2984 29880 2990
rect 29828 2926 29880 2932
rect 29644 2508 29696 2514
rect 29644 2450 29696 2456
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 30116 800 30144 2450
rect 30208 2446 30236 4966
rect 30300 4486 30328 6326
rect 30392 6322 30420 8230
rect 30576 8214 30696 8242
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30484 6662 30512 6734
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 30576 3890 30604 8214
rect 30760 7954 30788 8366
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30668 6866 30696 7822
rect 30852 7818 30880 8570
rect 30944 8090 30972 10610
rect 31036 9926 31064 11086
rect 31220 10198 31248 11562
rect 31208 10192 31260 10198
rect 31208 10134 31260 10140
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 30840 7812 30892 7818
rect 30840 7754 30892 7760
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30668 5234 30696 6802
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30654 5128 30710 5137
rect 30654 5063 30656 5072
rect 30708 5063 30710 5072
rect 30656 5034 30708 5040
rect 30760 4146 30788 7482
rect 30852 7324 30880 7754
rect 30944 7546 30972 7822
rect 31036 7818 31064 9522
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31128 8498 31156 9318
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 31024 7812 31076 7818
rect 31024 7754 31076 7760
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 30852 7296 31064 7324
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 30840 5568 30892 5574
rect 30840 5510 30892 5516
rect 30852 5234 30880 5510
rect 30944 5234 30972 6598
rect 31036 5710 31064 7296
rect 31128 6662 31156 7822
rect 31220 6866 31248 8026
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 31312 5302 31340 12786
rect 31588 12714 31616 14214
rect 31772 14006 31800 14214
rect 31760 14000 31812 14006
rect 31760 13942 31812 13948
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31576 12708 31628 12714
rect 31576 12650 31628 12656
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31404 12434 31432 12582
rect 31404 12406 31524 12434
rect 31496 12170 31524 12406
rect 31484 12164 31536 12170
rect 31484 12106 31536 12112
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31404 10266 31432 10678
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31404 8498 31432 10202
rect 31588 9586 31616 12650
rect 31680 12170 31708 13874
rect 31956 13394 31984 15642
rect 32140 15502 32168 15846
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32324 14822 32352 15302
rect 32508 14822 32536 16050
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 32312 14816 32364 14822
rect 32312 14758 32364 14764
rect 32496 14816 32548 14822
rect 32496 14758 32548 14764
rect 31944 13388 31996 13394
rect 31944 13330 31996 13336
rect 32324 12850 32352 14758
rect 32508 13530 32536 14758
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 33692 14068 33744 14074
rect 33692 14010 33744 14016
rect 32496 13524 32548 13530
rect 32496 13466 32548 13472
rect 32404 13320 32456 13326
rect 32404 13262 32456 13268
rect 32416 12850 32444 13262
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 32220 12640 32272 12646
rect 32220 12582 32272 12588
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31680 11830 31708 12106
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 31680 9722 31708 10610
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31772 9178 31800 9318
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 31404 8090 31432 8434
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7546 31432 7686
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31496 6934 31524 8434
rect 31576 7948 31628 7954
rect 31576 7890 31628 7896
rect 31588 7002 31616 7890
rect 31864 7478 31892 9454
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 31758 7032 31814 7041
rect 31576 6996 31628 7002
rect 31864 7002 31892 7414
rect 31758 6967 31814 6976
rect 31852 6996 31904 7002
rect 31576 6938 31628 6944
rect 31484 6928 31536 6934
rect 31484 6870 31536 6876
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 31116 5228 31168 5234
rect 31116 5170 31168 5176
rect 31128 4826 31156 5170
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31496 4622 31524 6870
rect 31772 5953 31800 6967
rect 31852 6938 31904 6944
rect 31956 6338 31984 10406
rect 32232 10282 32260 12582
rect 32324 10418 32352 12786
rect 32416 12434 32444 12786
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 32416 12406 32628 12434
rect 32600 12102 32628 12406
rect 32692 12238 32720 12582
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32324 10390 32536 10418
rect 32232 10254 32352 10282
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32036 9988 32088 9994
rect 32036 9930 32088 9936
rect 32048 9178 32076 9930
rect 32036 9172 32088 9178
rect 32036 9114 32088 9120
rect 32140 7886 32168 9998
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32232 9654 32260 9862
rect 32220 9648 32272 9654
rect 32220 9590 32272 9596
rect 32220 8968 32272 8974
rect 32220 8910 32272 8916
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32036 7744 32088 7750
rect 32036 7686 32088 7692
rect 32048 6390 32076 7686
rect 32232 6916 32260 8910
rect 32324 8906 32352 10254
rect 32508 10130 32536 10390
rect 32496 10124 32548 10130
rect 32496 10066 32548 10072
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 32416 9178 32444 9998
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 32312 8288 32364 8294
rect 32312 8230 32364 8236
rect 32324 7410 32352 8230
rect 32600 8022 32628 12038
rect 32692 11218 32720 12174
rect 33152 11778 33180 12786
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 33336 12238 33364 12718
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 33520 12594 33548 12650
rect 33428 12566 33548 12594
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32968 11750 33180 11778
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32784 10538 32812 11698
rect 32968 11694 32996 11750
rect 32956 11688 33008 11694
rect 32956 11630 33008 11636
rect 33152 10810 33180 11750
rect 33336 11558 33364 12174
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 33336 10742 33364 11494
rect 33324 10736 33376 10742
rect 33324 10678 33376 10684
rect 33428 10674 33456 12566
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 32772 10532 32824 10538
rect 32772 10474 32824 10480
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 33336 10248 33364 10542
rect 33416 10260 33468 10266
rect 33336 10220 33416 10248
rect 32968 10130 32996 10202
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 33232 10056 33284 10062
rect 33232 9998 33284 10004
rect 33060 9382 33088 9998
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 33048 9104 33100 9110
rect 33048 9046 33100 9052
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32692 8566 32720 8774
rect 33060 8650 33088 9046
rect 33152 8838 33180 9862
rect 33244 8974 33272 9998
rect 33336 9110 33364 10220
rect 33416 10202 33468 10208
rect 33520 10130 33548 11086
rect 33508 10124 33560 10130
rect 33508 10066 33560 10072
rect 33520 9722 33548 10066
rect 33600 9920 33652 9926
rect 33600 9862 33652 9868
rect 33508 9716 33560 9722
rect 33508 9658 33560 9664
rect 33324 9104 33376 9110
rect 33324 9046 33376 9052
rect 33416 9104 33468 9110
rect 33416 9046 33468 9052
rect 33232 8968 33284 8974
rect 33284 8916 33364 8922
rect 33232 8910 33364 8916
rect 33244 8894 33364 8910
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33060 8622 33180 8650
rect 32680 8560 32732 8566
rect 32680 8502 32732 8508
rect 33152 8498 33180 8622
rect 33232 8560 33284 8566
rect 33232 8502 33284 8508
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32496 7948 32548 7954
rect 32496 7890 32548 7896
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32416 7002 32444 7822
rect 32312 6996 32364 7002
rect 32312 6938 32364 6944
rect 32404 6996 32456 7002
rect 32404 6938 32456 6944
rect 32140 6888 32260 6916
rect 31864 6310 31984 6338
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 31758 5944 31814 5953
rect 31758 5879 31814 5888
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 31576 4480 31628 4486
rect 31576 4422 31628 4428
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30840 4140 30892 4146
rect 30892 4100 30972 4128
rect 30840 4082 30892 4088
rect 30760 4049 30788 4082
rect 30746 4040 30802 4049
rect 30746 3975 30802 3984
rect 30840 4004 30892 4010
rect 30840 3946 30892 3952
rect 30852 3890 30880 3946
rect 30576 3862 30880 3890
rect 30654 3496 30710 3505
rect 30654 3431 30656 3440
rect 30708 3431 30710 3440
rect 30656 3402 30708 3408
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 30852 3233 30880 3334
rect 30838 3224 30894 3233
rect 30472 3188 30524 3194
rect 30838 3159 30894 3168
rect 30472 3130 30524 3136
rect 30484 2650 30512 3130
rect 30944 3058 30972 4100
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30852 2961 30880 2994
rect 30838 2952 30894 2961
rect 30838 2887 30894 2896
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 31036 2446 31064 4422
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31116 4004 31168 4010
rect 31116 3946 31168 3952
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31128 3058 31156 3946
rect 31116 3052 31168 3058
rect 31116 2994 31168 3000
rect 31220 2990 31248 3946
rect 31312 3346 31340 4082
rect 31392 3936 31444 3942
rect 31392 3878 31444 3884
rect 31404 3466 31432 3878
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 31484 3460 31536 3466
rect 31484 3402 31536 3408
rect 31496 3346 31524 3402
rect 31312 3318 31524 3346
rect 31312 3058 31340 3318
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31588 2446 31616 4422
rect 31772 3233 31800 5646
rect 31864 5166 31892 6310
rect 31944 6180 31996 6186
rect 31944 6122 31996 6128
rect 31852 5160 31904 5166
rect 31852 5102 31904 5108
rect 31956 3505 31984 6122
rect 32140 5778 32168 6888
rect 32324 6848 32352 6938
rect 32232 6820 32352 6848
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 32232 4622 32260 6820
rect 32508 5166 32536 7890
rect 33048 7744 33100 7750
rect 33152 7732 33180 8434
rect 33244 7886 33272 8502
rect 33336 8362 33364 8894
rect 33324 8356 33376 8362
rect 33324 8298 33376 8304
rect 33428 8294 33456 9046
rect 33520 8974 33548 9658
rect 33612 9178 33640 9862
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33520 8566 33548 8910
rect 33612 8838 33640 9114
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 33508 8560 33560 8566
rect 33508 8502 33560 8508
rect 33612 8430 33640 8774
rect 33600 8424 33652 8430
rect 33600 8366 33652 8372
rect 33416 8288 33468 8294
rect 33416 8230 33468 8236
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33416 7812 33468 7818
rect 33416 7754 33468 7760
rect 33152 7704 33364 7732
rect 33048 7686 33100 7692
rect 33060 7478 33088 7686
rect 33048 7472 33100 7478
rect 33048 7414 33100 7420
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33152 6730 33180 6802
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33232 6724 33284 6730
rect 33232 6666 33284 6672
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32600 5574 32628 5714
rect 32692 5642 32720 6258
rect 32680 5636 32732 5642
rect 32680 5578 32732 5584
rect 32864 5636 32916 5642
rect 32864 5578 32916 5584
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32876 5098 32904 5578
rect 32864 5092 32916 5098
rect 32864 5034 32916 5040
rect 32220 4616 32272 4622
rect 32220 4558 32272 4564
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32140 4049 32168 4082
rect 32126 4040 32182 4049
rect 32126 3975 32182 3984
rect 32232 3534 32260 4558
rect 32312 4480 32364 4486
rect 32312 4422 32364 4428
rect 32324 4298 32352 4422
rect 32324 4270 32536 4298
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32324 3602 32352 4082
rect 32508 3942 32536 4270
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32312 3596 32364 3602
rect 32312 3538 32364 3544
rect 32220 3528 32272 3534
rect 31942 3496 31998 3505
rect 32220 3470 32272 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31942 3431 31998 3440
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 31758 3224 31814 3233
rect 31758 3159 31814 3168
rect 32324 2961 32352 3402
rect 32416 3058 32444 3470
rect 32600 3398 32628 4082
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32588 3392 32640 3398
rect 32588 3334 32640 3340
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32310 2952 32366 2961
rect 32310 2887 32366 2896
rect 32508 2774 32536 3130
rect 32692 3058 32720 3878
rect 32968 3602 32996 4014
rect 33060 3602 33088 6326
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 33152 4826 33180 6258
rect 33244 5370 33272 6666
rect 33232 5364 33284 5370
rect 33232 5306 33284 5312
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 32956 3596 33008 3602
rect 32956 3538 33008 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33152 3534 33180 4082
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 32680 3052 32732 3058
rect 32680 2994 32732 3000
rect 33152 2854 33180 3470
rect 33232 3460 33284 3466
rect 33336 3448 33364 7704
rect 33428 5710 33456 7754
rect 33600 7744 33652 7750
rect 33600 7686 33652 7692
rect 33612 7410 33640 7686
rect 33600 7404 33652 7410
rect 33600 7346 33652 7352
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33520 4593 33548 6598
rect 33704 6322 33732 14010
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 33876 12776 33928 12782
rect 33876 12718 33928 12724
rect 33888 11286 33916 12718
rect 33968 12640 34020 12646
rect 33968 12582 34020 12588
rect 33876 11280 33928 11286
rect 33876 11222 33928 11228
rect 33784 9988 33836 9994
rect 33784 9930 33836 9936
rect 33796 8906 33824 9930
rect 33888 9518 33916 11222
rect 33980 11150 34008 12582
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34152 11688 34204 11694
rect 34152 11630 34204 11636
rect 34164 11354 34192 11630
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 36268 11552 36320 11558
rect 36268 11494 36320 11500
rect 34152 11348 34204 11354
rect 34152 11290 34204 11296
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 34152 11144 34204 11150
rect 34152 11086 34204 11092
rect 34164 10538 34192 11086
rect 34244 10804 34296 10810
rect 34244 10746 34296 10752
rect 34152 10532 34204 10538
rect 34152 10474 34204 10480
rect 34152 10056 34204 10062
rect 34152 9998 34204 10004
rect 34060 9920 34112 9926
rect 34164 9897 34192 9998
rect 34060 9862 34112 9868
rect 34150 9888 34206 9897
rect 33876 9512 33928 9518
rect 33876 9454 33928 9460
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 33888 8922 33916 9318
rect 34072 9042 34100 9862
rect 34150 9823 34206 9832
rect 34256 9586 34284 10746
rect 34440 10674 34468 11494
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 34440 10062 34468 10610
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34428 10056 34480 10062
rect 34428 9998 34480 10004
rect 34624 9654 34652 10406
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 36280 10062 36308 11494
rect 36268 10056 36320 10062
rect 36268 9998 36320 10004
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 34612 9648 34664 9654
rect 34612 9590 34664 9596
rect 35636 9586 35664 9862
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 34612 9512 34664 9518
rect 34612 9454 34664 9460
rect 35440 9512 35492 9518
rect 35440 9454 35492 9460
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 34060 9036 34112 9042
rect 34060 8978 34112 8984
rect 33888 8906 34008 8922
rect 33784 8900 33836 8906
rect 33888 8900 34020 8906
rect 33888 8894 33968 8900
rect 33784 8842 33836 8848
rect 33968 8842 34020 8848
rect 34164 8566 34192 9318
rect 34532 8974 34560 9318
rect 34624 9178 34652 9454
rect 34796 9444 34848 9450
rect 34796 9386 34848 9392
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34440 8634 34468 8842
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34532 8498 34560 8910
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 33968 8356 34020 8362
rect 33968 8298 34020 8304
rect 33980 7206 34008 8298
rect 34060 7948 34112 7954
rect 34060 7890 34112 7896
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33692 6316 33744 6322
rect 33692 6258 33744 6264
rect 33690 5808 33746 5817
rect 33690 5743 33746 5752
rect 33704 5710 33732 5743
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33876 5568 33928 5574
rect 33876 5510 33928 5516
rect 33888 5234 33916 5510
rect 33980 5302 34008 7142
rect 33968 5296 34020 5302
rect 33968 5238 34020 5244
rect 33600 5228 33652 5234
rect 33600 5170 33652 5176
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 33612 4826 33640 5170
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 33506 4584 33562 4593
rect 33888 4554 33916 5170
rect 34072 5137 34100 7890
rect 34612 7880 34664 7886
rect 34612 7822 34664 7828
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34532 7313 34560 7686
rect 34518 7304 34574 7313
rect 34518 7239 34574 7248
rect 34624 7041 34652 7822
rect 34716 7410 34744 8910
rect 34808 8838 34836 9386
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34808 8498 34836 8774
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34610 7032 34666 7041
rect 34610 6967 34666 6976
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 5914 34284 6258
rect 34244 5908 34296 5914
rect 34244 5850 34296 5856
rect 34716 5778 34744 7346
rect 34808 6798 34836 8434
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 35360 7886 35388 8026
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35348 7540 35400 7546
rect 35348 7482 35400 7488
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 35256 6792 35308 6798
rect 35360 6746 35388 7482
rect 35452 6866 35480 9454
rect 35636 8362 35664 9522
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 35820 9178 35848 9318
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35624 8356 35676 8362
rect 35624 8298 35676 8304
rect 35532 8288 35584 8294
rect 35532 8230 35584 8236
rect 35544 7478 35572 8230
rect 35532 7472 35584 7478
rect 35532 7414 35584 7420
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 35308 6740 35388 6746
rect 35256 6734 35388 6740
rect 35072 6724 35124 6730
rect 35268 6718 35388 6734
rect 35072 6666 35124 6672
rect 34796 6452 34848 6458
rect 34796 6394 34848 6400
rect 34704 5772 34756 5778
rect 34704 5714 34756 5720
rect 34612 5704 34664 5710
rect 34610 5672 34612 5681
rect 34664 5672 34666 5681
rect 34610 5607 34666 5616
rect 34244 5568 34296 5574
rect 34244 5510 34296 5516
rect 34256 5370 34284 5510
rect 34244 5364 34296 5370
rect 34244 5306 34296 5312
rect 34716 5234 34744 5714
rect 34808 5302 34836 6394
rect 35084 6390 35112 6666
rect 35164 6452 35216 6458
rect 35164 6394 35216 6400
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 35176 6322 35204 6394
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35360 6254 35388 6718
rect 35636 6458 35664 8298
rect 35716 7744 35768 7750
rect 35716 7686 35768 7692
rect 35728 7002 35756 7686
rect 35716 6996 35768 7002
rect 35716 6938 35768 6944
rect 35820 6458 35848 8434
rect 36004 8430 36032 9522
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 35900 7200 35952 7206
rect 35900 7142 35952 7148
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35912 7002 35940 7142
rect 35900 6996 35952 7002
rect 35900 6938 35952 6944
rect 36004 6730 36032 7142
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 35900 6656 35952 6662
rect 35952 6604 36032 6610
rect 35900 6598 36032 6604
rect 35912 6582 36032 6598
rect 35624 6452 35676 6458
rect 35624 6394 35676 6400
rect 35808 6452 35860 6458
rect 35808 6394 35860 6400
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35716 6316 35768 6322
rect 35716 6258 35768 6264
rect 35348 6248 35400 6254
rect 35348 6190 35400 6196
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35636 5370 35664 6258
rect 35624 5364 35676 5370
rect 35624 5306 35676 5312
rect 34796 5296 34848 5302
rect 34796 5238 34848 5244
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 34058 5128 34114 5137
rect 34058 5063 34114 5072
rect 34520 5092 34572 5098
rect 33506 4519 33562 4528
rect 33876 4548 33928 4554
rect 33876 4490 33928 4496
rect 34072 4146 34100 5063
rect 34520 5034 34572 5040
rect 33508 4140 33560 4146
rect 33508 4082 33560 4088
rect 34060 4140 34112 4146
rect 34060 4082 34112 4088
rect 33520 3738 33548 4082
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33888 3738 33916 3878
rect 33508 3732 33560 3738
rect 33508 3674 33560 3680
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 33284 3420 33364 3448
rect 33232 3402 33284 3408
rect 34532 3398 34560 5034
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 33784 2984 33836 2990
rect 33784 2926 33836 2932
rect 33416 2916 33468 2922
rect 33416 2858 33468 2864
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 32416 2746 32536 2774
rect 31668 2576 31720 2582
rect 31668 2518 31720 2524
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30852 800 30880 2246
rect 31680 1170 31708 2518
rect 32416 1170 32444 2746
rect 32784 2514 32812 2790
rect 32772 2508 32824 2514
rect 32772 2450 32824 2456
rect 33428 2446 33456 2858
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33140 2304 33192 2310
rect 31588 1142 31708 1170
rect 32324 1142 32444 1170
rect 33060 2252 33140 2258
rect 33060 2246 33192 2252
rect 33060 2230 33180 2246
rect 31588 800 31616 1142
rect 32324 800 32352 1142
rect 33060 800 33088 2230
rect 33796 800 33824 2926
rect 34532 2650 34560 3130
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34624 2514 34652 3878
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 34716 2446 34744 3674
rect 34808 3534 34836 5238
rect 35440 5024 35492 5030
rect 35440 4966 35492 4972
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35070 4720 35126 4729
rect 35070 4655 35126 4664
rect 35084 4146 35112 4655
rect 35072 4140 35124 4146
rect 35072 4082 35124 4088
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 34808 3126 34836 3334
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34992 3058 35020 3538
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 34796 2916 34848 2922
rect 34796 2858 34848 2864
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 34808 1578 34836 2858
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34624 1550 34836 1578
rect 34624 800 34652 1550
rect 35360 800 35388 3878
rect 35452 2990 35480 4966
rect 35728 4622 35756 6258
rect 36004 6254 36032 6582
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 35808 5024 35860 5030
rect 35808 4966 35860 4972
rect 35820 4622 35848 4966
rect 35716 4616 35768 4622
rect 35716 4558 35768 4564
rect 35808 4616 35860 4622
rect 35808 4558 35860 4564
rect 35624 4480 35676 4486
rect 35624 4422 35676 4428
rect 35636 4214 35664 4422
rect 35624 4208 35676 4214
rect 35624 4150 35676 4156
rect 35636 3602 35664 4150
rect 35624 3596 35676 3602
rect 35624 3538 35676 3544
rect 35728 3534 35756 4558
rect 35912 4078 35940 5170
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35820 3126 35848 3334
rect 35808 3120 35860 3126
rect 35808 3062 35860 3068
rect 36004 3058 36032 6190
rect 36188 6186 36216 7822
rect 36268 6792 36320 6798
rect 36266 6760 36268 6769
rect 36728 6792 36780 6798
rect 36320 6760 36322 6769
rect 36728 6734 36780 6740
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 36266 6695 36322 6704
rect 36268 6656 36320 6662
rect 36268 6598 36320 6604
rect 36280 6390 36308 6598
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 36176 6180 36228 6186
rect 36176 6122 36228 6128
rect 36176 5908 36228 5914
rect 36096 5868 36176 5896
rect 36096 5642 36124 5868
rect 36176 5850 36228 5856
rect 36174 5672 36230 5681
rect 36084 5636 36136 5642
rect 36174 5607 36230 5616
rect 36084 5578 36136 5584
rect 36188 3534 36216 5607
rect 36280 4554 36308 6326
rect 36740 5817 36768 6734
rect 37188 6656 37240 6662
rect 37188 6598 37240 6604
rect 36726 5808 36782 5817
rect 36726 5743 36782 5752
rect 36728 5704 36780 5710
rect 36728 5646 36780 5652
rect 36452 4616 36504 4622
rect 36452 4558 36504 4564
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36268 4548 36320 4554
rect 36268 4490 36320 4496
rect 36464 3738 36492 4558
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 36096 800 36124 3334
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36188 2446 36216 2790
rect 36372 2650 36400 3130
rect 36556 2990 36584 4558
rect 36636 4140 36688 4146
rect 36636 4082 36688 4088
rect 36648 3670 36676 4082
rect 36636 3664 36688 3670
rect 36636 3606 36688 3612
rect 36636 3052 36688 3058
rect 36740 3040 36768 5646
rect 36912 5568 36964 5574
rect 36912 5510 36964 5516
rect 36924 4690 36952 5510
rect 37200 5302 37228 6598
rect 37188 5296 37240 5302
rect 37188 5238 37240 5244
rect 37384 4826 37412 6734
rect 37464 6112 37516 6118
rect 37464 6054 37516 6060
rect 37372 4820 37424 4826
rect 37372 4762 37424 4768
rect 37280 4752 37332 4758
rect 37476 4706 37504 6054
rect 37832 5840 37884 5846
rect 37832 5782 37884 5788
rect 37844 5234 37872 5782
rect 37832 5228 37884 5234
rect 37832 5170 37884 5176
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 39764 5024 39816 5030
rect 39764 4966 39816 4972
rect 37280 4694 37332 4700
rect 36912 4684 36964 4690
rect 36912 4626 36964 4632
rect 37292 3058 37320 4694
rect 37384 4678 37504 4706
rect 36688 3012 36768 3040
rect 37280 3052 37332 3058
rect 36636 2994 36688 3000
rect 37280 2994 37332 3000
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 36832 800 36860 2790
rect 37384 2446 37412 4678
rect 37844 4622 37872 4966
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37832 4480 37884 4486
rect 37832 4422 37884 4428
rect 39028 4480 39080 4486
rect 39028 4422 39080 4428
rect 37844 4146 37872 4422
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 38292 3936 38344 3942
rect 38292 3878 38344 3884
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37476 2650 37504 2926
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37568 800 37596 3334
rect 38304 800 38332 3878
rect 39040 800 39068 4422
rect 39776 800 39804 4966
rect 19720 734 19932 762
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3146 4392 3202 4448
rect 3054 3612 3056 3632
rect 3056 3612 3108 3632
rect 3108 3612 3110 3632
rect 3054 3576 3110 3612
rect 2686 3440 2742 3496
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 2226 2916 2282 2952
rect 2226 2896 2228 2916
rect 2228 2896 2280 2916
rect 2280 2896 2282 2916
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5538 5208 5594 5264
rect 4618 3884 4620 3904
rect 4620 3884 4672 3904
rect 4672 3884 4674 3904
rect 4618 3848 4674 3884
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4158 3168 4214 3224
rect 4434 3052 4490 3088
rect 4434 3032 4436 3052
rect 4436 3032 4488 3052
rect 4488 3032 4490 3052
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2352 4122 2408
rect 4894 3984 4950 4040
rect 5078 4256 5134 4312
rect 4802 3440 4858 3496
rect 4894 3304 4950 3360
rect 5354 4548 5410 4584
rect 5354 4528 5356 4548
rect 5356 4528 5408 4548
rect 5408 4528 5410 4548
rect 5262 4120 5318 4176
rect 5446 3576 5502 3632
rect 5814 4392 5870 4448
rect 5906 2216 5962 2272
rect 6274 4664 6330 4720
rect 6274 3712 6330 3768
rect 6734 4800 6790 4856
rect 6458 3712 6514 3768
rect 7378 4120 7434 4176
rect 7470 2760 7526 2816
rect 7838 3340 7840 3360
rect 7840 3340 7892 3360
rect 7892 3340 7894 3360
rect 7838 3304 7894 3340
rect 8206 2760 8262 2816
rect 8390 2488 8446 2544
rect 8942 7520 8998 7576
rect 10506 11056 10562 11112
rect 9494 5212 9550 5264
rect 9494 5208 9496 5212
rect 9496 5208 9548 5212
rect 9548 5208 9550 5212
rect 9862 5072 9918 5128
rect 10230 5072 10286 5128
rect 10138 4528 10194 4584
rect 9678 4140 9734 4176
rect 9678 4120 9680 4140
rect 9680 4120 9732 4140
rect 9732 4120 9734 4140
rect 8942 2352 8998 2408
rect 9494 3576 9550 3632
rect 9770 3576 9826 3632
rect 10046 3576 10102 3632
rect 10230 4120 10286 4176
rect 10690 3032 10746 3088
rect 13174 11076 13230 11112
rect 13174 11056 13176 11076
rect 13176 11056 13228 11076
rect 13228 11056 13230 11076
rect 11334 4256 11390 4312
rect 12254 3848 12310 3904
rect 16210 12280 16266 12336
rect 14830 12164 14886 12200
rect 14830 12144 14832 12164
rect 14832 12144 14884 12164
rect 14884 12144 14886 12164
rect 14922 8472 14978 8528
rect 13910 4664 13966 4720
rect 12530 3440 12586 3496
rect 13266 2488 13322 2544
rect 12806 2352 12862 2408
rect 13910 3712 13966 3768
rect 15290 5344 15346 5400
rect 14922 3984 14978 4040
rect 15014 3168 15070 3224
rect 15474 4800 15530 4856
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 17498 12164 17554 12200
rect 17498 12144 17500 12164
rect 17500 12144 17552 12164
rect 17552 12144 17554 12164
rect 17130 8472 17186 8528
rect 16854 5072 16910 5128
rect 18050 12300 18106 12336
rect 18050 12280 18052 12300
rect 18052 12280 18104 12300
rect 18104 12280 18106 12300
rect 18786 7520 18842 7576
rect 17038 2896 17094 2952
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19430 9016 19486 9072
rect 19706 9288 19762 9344
rect 20534 12164 20590 12200
rect 20534 12144 20536 12164
rect 20536 12144 20588 12164
rect 20588 12144 20590 12164
rect 20350 10532 20406 10568
rect 20350 10512 20352 10532
rect 20352 10512 20404 10532
rect 20404 10512 20406 10532
rect 20350 9288 20406 9344
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19890 7928 19946 7984
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20166 8064 20222 8120
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20902 5636 20958 5672
rect 20902 5616 20904 5636
rect 20904 5616 20956 5636
rect 20956 5616 20958 5636
rect 22098 9596 22100 9616
rect 22100 9596 22152 9616
rect 22152 9596 22154 9616
rect 22098 9560 22154 9596
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22742 9424 22798 9480
rect 22558 5772 22614 5808
rect 22558 5752 22560 5772
rect 22560 5752 22612 5772
rect 22612 5752 22614 5772
rect 22926 6432 22982 6488
rect 23938 10512 23994 10568
rect 23754 9560 23810 9616
rect 23570 9016 23626 9072
rect 23386 4548 23442 4584
rect 23386 4528 23388 4548
rect 23388 4528 23440 4548
rect 23440 4528 23442 4548
rect 24766 8084 24822 8120
rect 24766 8064 24768 8084
rect 24768 8064 24820 8084
rect 24820 8064 24822 8084
rect 25318 7948 25374 7984
rect 25318 7928 25320 7948
rect 25320 7928 25372 7948
rect 25372 7928 25374 7948
rect 25502 8608 25558 8664
rect 25594 8492 25650 8528
rect 25594 8472 25596 8492
rect 25596 8472 25648 8492
rect 25648 8472 25650 8492
rect 25410 5616 25466 5672
rect 25962 4140 26018 4176
rect 25962 4120 25964 4140
rect 25964 4120 26016 4140
rect 26016 4120 26018 4140
rect 26606 8608 26662 8664
rect 27526 8492 27582 8528
rect 27526 8472 27528 8492
rect 27528 8472 27580 8492
rect 27580 8472 27582 8492
rect 27342 5888 27398 5944
rect 27342 3460 27398 3496
rect 27342 3440 27344 3460
rect 27344 3440 27396 3460
rect 27396 3440 27398 3460
rect 27986 6724 28042 6760
rect 27986 6704 27988 6724
rect 27988 6704 28040 6724
rect 28040 6704 28042 6724
rect 28630 12164 28686 12200
rect 28630 12144 28632 12164
rect 28632 12144 28684 12164
rect 28684 12144 28686 12164
rect 28446 8200 28502 8256
rect 28722 9444 28778 9480
rect 28722 9424 28724 9444
rect 28724 9424 28776 9444
rect 28776 9424 28778 9444
rect 28814 8200 28870 8256
rect 28814 8064 28870 8120
rect 28998 7928 29054 7984
rect 28262 6432 28318 6488
rect 28170 5480 28226 5536
rect 28170 3476 28172 3496
rect 28172 3476 28224 3496
rect 28224 3476 28226 3496
rect 28170 3440 28226 3476
rect 28170 2896 28226 2952
rect 28906 4140 28962 4176
rect 28906 4120 28908 4140
rect 28908 4120 28960 4140
rect 28960 4120 28962 4140
rect 30378 9832 30434 9888
rect 29366 4664 29422 4720
rect 30654 5092 30710 5128
rect 30654 5072 30656 5092
rect 30656 5072 30708 5092
rect 30708 5072 30710 5092
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 31758 6976 31814 7032
rect 31758 5888 31814 5944
rect 30746 3984 30802 4040
rect 30654 3460 30710 3496
rect 30654 3440 30656 3460
rect 30656 3440 30708 3460
rect 30708 3440 30710 3460
rect 30838 3168 30894 3224
rect 30838 2896 30894 2952
rect 32126 3984 32182 4040
rect 31942 3440 31998 3496
rect 31758 3168 31814 3224
rect 32310 2896 32366 2952
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34150 9832 34206 9888
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 33690 5752 33746 5808
rect 33506 4528 33562 4584
rect 34518 7248 34574 7304
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34610 6976 34666 7032
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34610 5652 34612 5672
rect 34612 5652 34664 5672
rect 34664 5652 34666 5672
rect 34610 5616 34666 5652
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34058 5072 34114 5128
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35070 4664 35126 4720
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36266 6740 36268 6760
rect 36268 6740 36320 6760
rect 36320 6740 36322 6760
rect 36266 6704 36322 6740
rect 36174 5616 36230 5672
rect 36726 5752 36782 5808
<< metal3 >>
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25032 800 25152
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 16205 12338 16271 12341
rect 18045 12338 18111 12341
rect 16205 12336 18111 12338
rect 16205 12280 16210 12336
rect 16266 12280 18050 12336
rect 18106 12280 18111 12336
rect 16205 12278 18111 12280
rect 16205 12275 16271 12278
rect 18045 12275 18111 12278
rect 14825 12202 14891 12205
rect 17493 12202 17559 12205
rect 14825 12200 17559 12202
rect 14825 12144 14830 12200
rect 14886 12144 17498 12200
rect 17554 12144 17559 12200
rect 14825 12142 17559 12144
rect 14825 12139 14891 12142
rect 17493 12139 17559 12142
rect 20529 12202 20595 12205
rect 28625 12202 28691 12205
rect 20529 12200 28691 12202
rect 20529 12144 20534 12200
rect 20590 12144 28630 12200
rect 28686 12144 28691 12200
rect 20529 12142 28691 12144
rect 20529 12139 20595 12142
rect 28625 12139 28691 12142
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 10501 11114 10567 11117
rect 13169 11114 13235 11117
rect 10501 11112 13235 11114
rect 10501 11056 10506 11112
rect 10562 11056 13174 11112
rect 13230 11056 13235 11112
rect 10501 11054 13235 11056
rect 10501 11051 10567 11054
rect 13169 11051 13235 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 20345 10570 20411 10573
rect 23933 10570 23999 10573
rect 20345 10568 23999 10570
rect 20345 10512 20350 10568
rect 20406 10512 23938 10568
rect 23994 10512 23999 10568
rect 20345 10510 23999 10512
rect 20345 10507 20411 10510
rect 23933 10507 23999 10510
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 30373 9890 30439 9893
rect 34145 9890 34211 9893
rect 30373 9888 34211 9890
rect 30373 9832 30378 9888
rect 30434 9832 34150 9888
rect 34206 9832 34211 9888
rect 30373 9830 34211 9832
rect 30373 9827 30439 9830
rect 34145 9827 34211 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 22093 9618 22159 9621
rect 23749 9618 23815 9621
rect 22093 9616 23815 9618
rect 22093 9560 22098 9616
rect 22154 9560 23754 9616
rect 23810 9560 23815 9616
rect 22093 9558 23815 9560
rect 22093 9555 22159 9558
rect 23749 9555 23815 9558
rect 22737 9482 22803 9485
rect 28717 9482 28783 9485
rect 22737 9480 28783 9482
rect 22737 9424 22742 9480
rect 22798 9424 28722 9480
rect 28778 9424 28783 9480
rect 22737 9422 28783 9424
rect 22737 9419 22803 9422
rect 28717 9419 28783 9422
rect 19701 9346 19767 9349
rect 20345 9346 20411 9349
rect 19701 9344 20411 9346
rect 19701 9288 19706 9344
rect 19762 9288 20350 9344
rect 20406 9288 20411 9344
rect 19701 9286 20411 9288
rect 19701 9283 19767 9286
rect 20345 9283 20411 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 19425 9074 19491 9077
rect 23565 9074 23631 9077
rect 19425 9072 23631 9074
rect 19425 9016 19430 9072
rect 19486 9016 23570 9072
rect 23626 9016 23631 9072
rect 19425 9014 23631 9016
rect 19425 9011 19491 9014
rect 23565 9011 23631 9014
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 25497 8666 25563 8669
rect 26601 8666 26667 8669
rect 25497 8664 26667 8666
rect 25497 8608 25502 8664
rect 25558 8608 26606 8664
rect 26662 8608 26667 8664
rect 25497 8606 26667 8608
rect 25497 8603 25563 8606
rect 26601 8603 26667 8606
rect 14917 8530 14983 8533
rect 17125 8530 17191 8533
rect 14917 8528 17191 8530
rect 14917 8472 14922 8528
rect 14978 8472 17130 8528
rect 17186 8472 17191 8528
rect 14917 8470 17191 8472
rect 14917 8467 14983 8470
rect 17125 8467 17191 8470
rect 25589 8530 25655 8533
rect 27521 8530 27587 8533
rect 25589 8528 27587 8530
rect 25589 8472 25594 8528
rect 25650 8472 27526 8528
rect 27582 8472 27587 8528
rect 25589 8470 27587 8472
rect 25589 8467 25655 8470
rect 27521 8467 27587 8470
rect 28441 8258 28507 8261
rect 28809 8258 28875 8261
rect 28441 8256 28875 8258
rect 28441 8200 28446 8256
rect 28502 8200 28814 8256
rect 28870 8200 28875 8256
rect 28441 8198 28875 8200
rect 28441 8195 28507 8198
rect 28809 8195 28875 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 20161 8122 20227 8125
rect 24761 8122 24827 8125
rect 28809 8122 28875 8125
rect 20161 8120 28875 8122
rect 20161 8064 20166 8120
rect 20222 8064 24766 8120
rect 24822 8064 28814 8120
rect 28870 8064 28875 8120
rect 20161 8062 28875 8064
rect 20161 8059 20227 8062
rect 24761 8059 24827 8062
rect 28809 8059 28875 8062
rect 19885 7986 19951 7989
rect 25313 7986 25379 7989
rect 28993 7986 29059 7989
rect 19885 7984 29059 7986
rect 19885 7928 19890 7984
rect 19946 7928 25318 7984
rect 25374 7928 28998 7984
rect 29054 7928 29059 7984
rect 19885 7926 29059 7928
rect 19885 7923 19951 7926
rect 25313 7923 25379 7926
rect 28993 7923 29059 7926
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 8937 7578 9003 7581
rect 18781 7578 18847 7581
rect 8937 7576 18847 7578
rect 8937 7520 8942 7576
rect 8998 7520 18786 7576
rect 18842 7520 18847 7576
rect 8937 7518 18847 7520
rect 8937 7515 9003 7518
rect 18781 7515 18847 7518
rect 30414 7244 30420 7308
rect 30484 7306 30490 7308
rect 34513 7306 34579 7309
rect 30484 7304 34579 7306
rect 30484 7248 34518 7304
rect 34574 7248 34579 7304
rect 30484 7246 34579 7248
rect 30484 7244 30490 7246
rect 34513 7243 34579 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 31753 7034 31819 7037
rect 34605 7034 34671 7037
rect 31753 7032 34671 7034
rect 31753 6976 31758 7032
rect 31814 6976 34610 7032
rect 34666 6976 34671 7032
rect 31753 6974 34671 6976
rect 31753 6971 31819 6974
rect 34605 6971 34671 6974
rect 27981 6762 28047 6765
rect 36261 6762 36327 6765
rect 27981 6760 36327 6762
rect 27981 6704 27986 6760
rect 28042 6704 36266 6760
rect 36322 6704 36327 6760
rect 27981 6702 36327 6704
rect 27981 6699 28047 6702
rect 36261 6699 36327 6702
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 22921 6490 22987 6493
rect 28257 6490 28323 6493
rect 22921 6488 28323 6490
rect 22921 6432 22926 6488
rect 22982 6432 28262 6488
rect 28318 6432 28323 6488
rect 22921 6430 28323 6432
rect 22921 6427 22987 6430
rect 28257 6427 28323 6430
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 27337 5946 27403 5949
rect 31753 5946 31819 5949
rect 27337 5944 31819 5946
rect 27337 5888 27342 5944
rect 27398 5888 31758 5944
rect 31814 5888 31819 5944
rect 27337 5886 31819 5888
rect 27337 5883 27403 5886
rect 31753 5883 31819 5886
rect 22553 5810 22619 5813
rect 33685 5810 33751 5813
rect 36721 5810 36787 5813
rect 22553 5808 36787 5810
rect 22553 5752 22558 5808
rect 22614 5752 33690 5808
rect 33746 5752 36726 5808
rect 36782 5752 36787 5808
rect 22553 5750 36787 5752
rect 22553 5747 22619 5750
rect 33685 5747 33751 5750
rect 36721 5747 36787 5750
rect 20897 5674 20963 5677
rect 25405 5674 25471 5677
rect 20897 5672 25471 5674
rect 20897 5616 20902 5672
rect 20958 5616 25410 5672
rect 25466 5616 25471 5672
rect 20897 5614 25471 5616
rect 20897 5611 20963 5614
rect 25405 5611 25471 5614
rect 34605 5674 34671 5677
rect 36169 5674 36235 5677
rect 34605 5672 36235 5674
rect 34605 5616 34610 5672
rect 34666 5616 36174 5672
rect 36230 5616 36235 5672
rect 34605 5614 36235 5616
rect 34605 5611 34671 5614
rect 36169 5611 36235 5614
rect 28165 5538 28231 5541
rect 30414 5538 30420 5540
rect 28165 5536 30420 5538
rect 28165 5480 28170 5536
rect 28226 5480 30420 5536
rect 28165 5478 30420 5480
rect 28165 5475 28231 5478
rect 30414 5476 30420 5478
rect 30484 5476 30490 5540
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 4654 5340 4660 5404
rect 4724 5402 4730 5404
rect 15285 5402 15351 5405
rect 4724 5400 15351 5402
rect 4724 5344 15290 5400
rect 15346 5344 15351 5400
rect 4724 5342 15351 5344
rect 4724 5340 4730 5342
rect 15285 5339 15351 5342
rect 5533 5266 5599 5269
rect 9489 5266 9555 5269
rect 5533 5264 9555 5266
rect 5533 5208 5538 5264
rect 5594 5208 9494 5264
rect 9550 5208 9555 5264
rect 5533 5206 9555 5208
rect 5533 5203 5599 5206
rect 9489 5203 9555 5206
rect 9857 5132 9923 5133
rect 9806 5130 9812 5132
rect 9766 5070 9812 5130
rect 9876 5128 9923 5132
rect 9918 5072 9923 5128
rect 9806 5068 9812 5070
rect 9876 5068 9923 5072
rect 9857 5067 9923 5068
rect 10225 5130 10291 5133
rect 16849 5130 16915 5133
rect 10225 5128 16915 5130
rect 10225 5072 10230 5128
rect 10286 5072 16854 5128
rect 16910 5072 16915 5128
rect 10225 5070 16915 5072
rect 10225 5067 10291 5070
rect 16849 5067 16915 5070
rect 30649 5130 30715 5133
rect 34053 5130 34119 5133
rect 30649 5128 34119 5130
rect 30649 5072 30654 5128
rect 30710 5072 34058 5128
rect 34114 5072 34119 5128
rect 30649 5070 34119 5072
rect 30649 5067 30715 5070
rect 34053 5067 34119 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 6729 4858 6795 4861
rect 15469 4858 15535 4861
rect 6729 4856 15535 4858
rect 6729 4800 6734 4856
rect 6790 4800 15474 4856
rect 15530 4800 15535 4856
rect 6729 4798 15535 4800
rect 6729 4795 6795 4798
rect 15469 4795 15535 4798
rect 6269 4722 6335 4725
rect 13905 4722 13971 4725
rect 6269 4720 13971 4722
rect 6269 4664 6274 4720
rect 6330 4664 13910 4720
rect 13966 4664 13971 4720
rect 6269 4662 13971 4664
rect 6269 4659 6335 4662
rect 13905 4659 13971 4662
rect 29361 4722 29427 4725
rect 35065 4722 35131 4725
rect 29361 4720 35131 4722
rect 29361 4664 29366 4720
rect 29422 4664 35070 4720
rect 35126 4664 35131 4720
rect 29361 4662 35131 4664
rect 29361 4659 29427 4662
rect 35065 4659 35131 4662
rect 5349 4586 5415 4589
rect 10133 4586 10199 4589
rect 5349 4584 10199 4586
rect 5349 4528 5354 4584
rect 5410 4528 10138 4584
rect 10194 4528 10199 4584
rect 5349 4526 10199 4528
rect 5349 4523 5415 4526
rect 10133 4523 10199 4526
rect 23381 4586 23447 4589
rect 33501 4586 33567 4589
rect 23381 4584 33567 4586
rect 23381 4528 23386 4584
rect 23442 4528 33506 4584
rect 33562 4528 33567 4584
rect 23381 4526 33567 4528
rect 23381 4523 23447 4526
rect 33501 4523 33567 4526
rect 3141 4450 3207 4453
rect 5809 4450 5875 4453
rect 3141 4448 5875 4450
rect 3141 4392 3146 4448
rect 3202 4392 5814 4448
rect 5870 4392 5875 4448
rect 3141 4390 5875 4392
rect 3141 4387 3207 4390
rect 5809 4387 5875 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 5073 4314 5139 4317
rect 11329 4314 11395 4317
rect 5073 4312 11395 4314
rect 5073 4256 5078 4312
rect 5134 4256 11334 4312
rect 11390 4256 11395 4312
rect 5073 4254 11395 4256
rect 5073 4251 5139 4254
rect 11329 4251 11395 4254
rect 5257 4178 5323 4181
rect 7373 4178 7439 4181
rect 5257 4176 7439 4178
rect 5257 4120 5262 4176
rect 5318 4120 7378 4176
rect 7434 4120 7439 4176
rect 5257 4118 7439 4120
rect 5257 4115 5323 4118
rect 7373 4115 7439 4118
rect 9673 4178 9739 4181
rect 10225 4178 10291 4181
rect 9673 4176 10291 4178
rect 9673 4120 9678 4176
rect 9734 4120 10230 4176
rect 10286 4120 10291 4176
rect 9673 4118 10291 4120
rect 9673 4115 9739 4118
rect 10225 4115 10291 4118
rect 25957 4178 26023 4181
rect 28901 4178 28967 4181
rect 25957 4176 28967 4178
rect 25957 4120 25962 4176
rect 26018 4120 28906 4176
rect 28962 4120 28967 4176
rect 25957 4118 28967 4120
rect 25957 4115 26023 4118
rect 28901 4115 28967 4118
rect 4889 4042 4955 4045
rect 14917 4042 14983 4045
rect 4889 4040 14983 4042
rect 4889 3984 4894 4040
rect 4950 3984 14922 4040
rect 14978 3984 14983 4040
rect 4889 3982 14983 3984
rect 4889 3979 4955 3982
rect 14917 3979 14983 3982
rect 30741 4042 30807 4045
rect 32121 4042 32187 4045
rect 30741 4040 32187 4042
rect 30741 3984 30746 4040
rect 30802 3984 32126 4040
rect 32182 3984 32187 4040
rect 30741 3982 32187 3984
rect 30741 3979 30807 3982
rect 32121 3979 32187 3982
rect 4613 3906 4679 3909
rect 12249 3906 12315 3909
rect 4613 3904 12315 3906
rect 4613 3848 4618 3904
rect 4674 3848 12254 3904
rect 12310 3848 12315 3904
rect 4613 3846 12315 3848
rect 4613 3843 4679 3846
rect 12249 3843 12315 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 6269 3770 6335 3773
rect 5214 3768 6335 3770
rect 5214 3712 6274 3768
rect 6330 3712 6335 3768
rect 5214 3710 6335 3712
rect 3049 3634 3115 3637
rect 5214 3634 5274 3710
rect 6269 3707 6335 3710
rect 6453 3770 6519 3773
rect 13905 3770 13971 3773
rect 6453 3768 13971 3770
rect 6453 3712 6458 3768
rect 6514 3712 13910 3768
rect 13966 3712 13971 3768
rect 6453 3710 13971 3712
rect 6453 3707 6519 3710
rect 13905 3707 13971 3710
rect 3049 3632 5274 3634
rect 3049 3576 3054 3632
rect 3110 3576 5274 3632
rect 3049 3574 5274 3576
rect 5441 3634 5507 3637
rect 9489 3634 9555 3637
rect 9765 3636 9831 3637
rect 9765 3634 9812 3636
rect 5441 3632 9555 3634
rect 5441 3576 5446 3632
rect 5502 3576 9494 3632
rect 9550 3576 9555 3632
rect 5441 3574 9555 3576
rect 9720 3632 9812 3634
rect 9876 3634 9882 3636
rect 10041 3634 10107 3637
rect 9876 3632 10107 3634
rect 9720 3576 9770 3632
rect 9876 3576 10046 3632
rect 10102 3576 10107 3632
rect 9720 3574 9812 3576
rect 3049 3571 3115 3574
rect 5441 3571 5507 3574
rect 9489 3571 9555 3574
rect 9765 3572 9812 3574
rect 9876 3574 10107 3576
rect 9876 3572 9882 3574
rect 9765 3571 9831 3572
rect 10041 3571 10107 3574
rect 2681 3498 2747 3501
rect 4654 3498 4660 3500
rect 2681 3496 4660 3498
rect 2681 3440 2686 3496
rect 2742 3440 4660 3496
rect 2681 3438 4660 3440
rect 2681 3435 2747 3438
rect 4654 3436 4660 3438
rect 4724 3436 4730 3500
rect 4797 3498 4863 3501
rect 12525 3498 12591 3501
rect 4797 3496 12591 3498
rect 4797 3440 4802 3496
rect 4858 3440 12530 3496
rect 12586 3440 12591 3496
rect 4797 3438 12591 3440
rect 4797 3435 4863 3438
rect 12525 3435 12591 3438
rect 27337 3498 27403 3501
rect 28165 3498 28231 3501
rect 27337 3496 28231 3498
rect 27337 3440 27342 3496
rect 27398 3440 28170 3496
rect 28226 3440 28231 3496
rect 27337 3438 28231 3440
rect 27337 3435 27403 3438
rect 28165 3435 28231 3438
rect 30649 3498 30715 3501
rect 31937 3498 32003 3501
rect 30649 3496 32003 3498
rect 30649 3440 30654 3496
rect 30710 3440 31942 3496
rect 31998 3440 32003 3496
rect 30649 3438 32003 3440
rect 30649 3435 30715 3438
rect 31937 3435 32003 3438
rect 4889 3362 4955 3365
rect 7833 3362 7899 3365
rect 4889 3360 7899 3362
rect 4889 3304 4894 3360
rect 4950 3304 7838 3360
rect 7894 3304 7899 3360
rect 4889 3302 7899 3304
rect 4889 3299 4955 3302
rect 7833 3299 7899 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4153 3226 4219 3229
rect 15009 3226 15075 3229
rect 4153 3224 15075 3226
rect 4153 3168 4158 3224
rect 4214 3168 15014 3224
rect 15070 3168 15075 3224
rect 4153 3166 15075 3168
rect 4153 3163 4219 3166
rect 15009 3163 15075 3166
rect 30833 3226 30899 3229
rect 31753 3226 31819 3229
rect 30833 3224 31819 3226
rect 30833 3168 30838 3224
rect 30894 3168 31758 3224
rect 31814 3168 31819 3224
rect 30833 3166 31819 3168
rect 30833 3163 30899 3166
rect 31753 3163 31819 3166
rect 4429 3090 4495 3093
rect 10685 3090 10751 3093
rect 4429 3088 10751 3090
rect 4429 3032 4434 3088
rect 4490 3032 10690 3088
rect 10746 3032 10751 3088
rect 4429 3030 10751 3032
rect 4429 3027 4495 3030
rect 10685 3027 10751 3030
rect 2221 2954 2287 2957
rect 17033 2954 17099 2957
rect 2221 2952 17099 2954
rect 2221 2896 2226 2952
rect 2282 2896 17038 2952
rect 17094 2896 17099 2952
rect 2221 2894 17099 2896
rect 2221 2891 2287 2894
rect 17033 2891 17099 2894
rect 28165 2954 28231 2957
rect 30833 2954 30899 2957
rect 32305 2954 32371 2957
rect 28165 2952 32371 2954
rect 28165 2896 28170 2952
rect 28226 2896 30838 2952
rect 30894 2896 32310 2952
rect 32366 2896 32371 2952
rect 28165 2894 32371 2896
rect 28165 2891 28231 2894
rect 30833 2891 30899 2894
rect 32305 2891 32371 2894
rect 7465 2818 7531 2821
rect 8201 2818 8267 2821
rect 7465 2816 8267 2818
rect 7465 2760 7470 2816
rect 7526 2760 8206 2816
rect 8262 2760 8267 2816
rect 7465 2758 8267 2760
rect 7465 2755 7531 2758
rect 8201 2755 8267 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 8385 2546 8451 2549
rect 13261 2546 13327 2549
rect 8385 2544 13327 2546
rect 8385 2488 8390 2544
rect 8446 2488 13266 2544
rect 13322 2488 13327 2544
rect 8385 2486 13327 2488
rect 8385 2483 8451 2486
rect 13261 2483 13327 2486
rect 4061 2410 4127 2413
rect 8937 2410 9003 2413
rect 12801 2410 12867 2413
rect 4061 2408 9003 2410
rect 4061 2352 4066 2408
rect 4122 2352 8942 2408
rect 8998 2352 9003 2408
rect 4061 2350 9003 2352
rect 4061 2347 4127 2350
rect 8937 2347 9003 2350
rect 12390 2408 12867 2410
rect 12390 2352 12806 2408
rect 12862 2352 12867 2408
rect 12390 2350 12867 2352
rect 5901 2274 5967 2277
rect 12390 2274 12450 2350
rect 12801 2347 12867 2350
rect 5901 2272 12450 2274
rect 5901 2216 5906 2272
rect 5962 2216 12450 2272
rect 5901 2214 12450 2216
rect 5901 2211 5967 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 30420 7244 30484 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 30420 5476 30484 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4660 5340 4724 5404
rect 9812 5128 9876 5132
rect 9812 5072 9862 5128
rect 9862 5072 9876 5128
rect 9812 5068 9876 5072
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 9812 3632 9876 3636
rect 9812 3576 9826 3632
rect 9826 3576 9876 3632
rect 9812 3572 9876 3576
rect 4660 3436 4724 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 30419 7308 30485 7309
rect 30419 7244 30420 7308
rect 30484 7244 30485 7308
rect 30419 7243 30485 7244
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 30422 5541 30482 7243
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 30419 5540 30485 5541
rect 30419 5476 30420 5540
rect 30484 5476 30485 5540
rect 30419 5475 30485 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 4659 5404 4725 5405
rect 4659 5340 4660 5404
rect 4724 5340 4725 5404
rect 4659 5339 4725 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4662 3501 4722 5339
rect 9811 5132 9877 5133
rect 9811 5068 9812 5132
rect 9876 5068 9877 5132
rect 9811 5067 9877 5068
rect 9814 3637 9874 5067
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 9811 3636 9877 3637
rect 9811 3572 9812 3636
rect 9876 3572 9877 3636
rect 9811 3571 9877 3572
rect 4659 3500 4725 3501
rect 4659 3436 4660 3500
rect 4724 3436 4725 3500
rect 4659 3435 4725 3436
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1644511149
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60
timestamp 1644511149
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1644511149
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96
timestamp 1644511149
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1644511149
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1644511149
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1644511149
transform 1 0 14720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1644511149
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1644511149
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1644511149
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1644511149
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_341
timestamp 1644511149
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1644511149
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_397
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1644511149
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_84
timestamp 1644511149
transform 1 0 8832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1644511149
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_201
timestamp 1644511149
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1644511149
transform 1 0 20792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_235
timestamp 1644511149
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_298
timestamp 1644511149
transform 1 0 28520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_307
timestamp 1644511149
transform 1 0 29348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_315
timestamp 1644511149
transform 1 0 30084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1644511149
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1644511149
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1644511149
transform 1 0 35328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_381
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1644511149
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1644511149
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1644511149
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1644511149
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_280
timestamp 1644511149
transform 1 0 26864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_314
timestamp 1644511149
transform 1 0 29992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1644511149
transform 1 0 32200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_351
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1644511149
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_379
timestamp 1644511149
transform 1 0 35972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_387
timestamp 1644511149
transform 1 0 36708 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1644511149
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_31
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_82
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1644511149
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_141
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_176
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1644511149
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1644511149
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_234
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_251
timestamp 1644511149
transform 1 0 24196 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1644511149
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1644511149
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_295
timestamp 1644511149
transform 1 0 28244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_299
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_314
timestamp 1644511149
transform 1 0 29992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_320
timestamp 1644511149
transform 1 0 30544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_346
timestamp 1644511149
transform 1 0 32936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_353
timestamp 1644511149
transform 1 0 33580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_360
timestamp 1644511149
transform 1 0 34224 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_366
timestamp 1644511149
transform 1 0 34776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_372
timestamp 1644511149
transform 1 0 35328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1644511149
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_6 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp 1644511149
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1644511149
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1644511149
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1644511149
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1644511149
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1644511149
transform 1 0 10764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_114
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_146
timestamp 1644511149
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1644511149
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1644511149
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_171
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1644511149
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1644511149
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_222
timestamp 1644511149
transform 1 0 21528 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_230
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1644511149
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1644511149
transform 1 0 26312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_281
timestamp 1644511149
transform 1 0 26956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1644511149
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_312
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_319
timestamp 1644511149
transform 1 0 30452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_326
timestamp 1644511149
transform 1 0 31096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_337
timestamp 1644511149
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1644511149
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1644511149
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_371
timestamp 1644511149
transform 1 0 35236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_378
timestamp 1644511149
transform 1 0 35880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_385
timestamp 1644511149
transform 1 0 36524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_391
timestamp 1644511149
transform 1 0 37076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1644511149
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1644511149
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1644511149
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1644511149
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1644511149
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1644511149
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1644511149
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_186
timestamp 1644511149
transform 1 0 18216 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_202
timestamp 1644511149
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_206
timestamp 1644511149
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1644511149
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_231
timestamp 1644511149
transform 1 0 22356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_246
timestamp 1644511149
transform 1 0 23736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_254
timestamp 1644511149
transform 1 0 24472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_262
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_270
timestamp 1644511149
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1644511149
transform 1 0 28704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_307
timestamp 1644511149
transform 1 0 29348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_315
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1644511149
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_341
timestamp 1644511149
transform 1 0 32476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_355
timestamp 1644511149
transform 1 0 33764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1644511149
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1644511149
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1644511149
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1644511149
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1644511149
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_182
timestamp 1644511149
transform 1 0 17848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1644511149
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_227
timestamp 1644511149
transform 1 0 21988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1644511149
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_272
timestamp 1644511149
transform 1 0 26128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_292
timestamp 1644511149
transform 1 0 27968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1644511149
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp 1644511149
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_335
timestamp 1644511149
transform 1 0 31924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_348
timestamp 1644511149
transform 1 0 33120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_355
timestamp 1644511149
transform 1 0 33764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1644511149
transform 1 0 36156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_388
timestamp 1644511149
transform 1 0 36800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1644511149
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_402
timestamp 1644511149
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1644511149
transform 1 0 38456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1644511149
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_60
timestamp 1644511149
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1644511149
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1644511149
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1644511149
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1644511149
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1644511149
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1644511149
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_175
timestamp 1644511149
transform 1 0 17204 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_182
timestamp 1644511149
transform 1 0 17848 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_204
timestamp 1644511149
transform 1 0 19872 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_229
timestamp 1644511149
transform 1 0 22172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_269
timestamp 1644511149
transform 1 0 25852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_288
timestamp 1644511149
transform 1 0 27600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_299
timestamp 1644511149
transform 1 0 28612 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_303
timestamp 1644511149
transform 1 0 28980 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1644511149
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_327
timestamp 1644511149
transform 1 0 31188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1644511149
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_357
timestamp 1644511149
transform 1 0 33948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_366
timestamp 1644511149
transform 1 0 34776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_377
timestamp 1644511149
transform 1 0 35788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1644511149
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1644511149
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_70
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_90
timestamp 1644511149
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_104
timestamp 1644511149
transform 1 0 10672 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_110
timestamp 1644511149
transform 1 0 11224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1644511149
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1644511149
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1644511149
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_160
timestamp 1644511149
transform 1 0 15824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_172
timestamp 1644511149
transform 1 0 16928 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_180
timestamp 1644511149
transform 1 0 17664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1644511149
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1644511149
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1644511149
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1644511149
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1644511149
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_271
timestamp 1644511149
transform 1 0 26036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_275
timestamp 1644511149
transform 1 0 26404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_282
timestamp 1644511149
transform 1 0 27048 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_293
timestamp 1644511149
transform 1 0 28060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_320
timestamp 1644511149
transform 1 0 30544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1644511149
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_348
timestamp 1644511149
transform 1 0 33120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1644511149
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_374
timestamp 1644511149
transform 1 0 35512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_381
timestamp 1644511149
transform 1 0 36156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1644511149
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_66
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_88
timestamp 1644511149
transform 1 0 9200 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1644511149
transform 1 0 9752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_124
timestamp 1644511149
transform 1 0 12512 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_130
timestamp 1644511149
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1644511149
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1644511149
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1644511149
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1644511149
transform 1 0 18308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_191
timestamp 1644511149
transform 1 0 18676 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_204
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_211
timestamp 1644511149
transform 1 0 20516 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_245
timestamp 1644511149
transform 1 0 23644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_253
timestamp 1644511149
transform 1 0 24380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_271
timestamp 1644511149
transform 1 0 26036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_298
timestamp 1644511149
transform 1 0 28520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_306
timestamp 1644511149
transform 1 0 29256 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1644511149
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_341
timestamp 1644511149
transform 1 0 32476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1644511149
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_364
timestamp 1644511149
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_381
timestamp 1644511149
transform 1 0 36156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1644511149
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1644511149
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_104
timestamp 1644511149
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1644511149
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1644511149
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1644511149
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp 1644511149
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_210
timestamp 1644511149
transform 1 0 20424 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1644511149
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_228
timestamp 1644511149
transform 1 0 22080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_257
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_278
timestamp 1644511149
transform 1 0 26680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1644511149
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1644511149
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_341
timestamp 1644511149
transform 1 0 32476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_349
timestamp 1644511149
transform 1 0 33212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1644511149
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_368
timestamp 1644511149
transform 1 0 34960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_375
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_382
timestamp 1644511149
transform 1 0 36248 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_394
timestamp 1644511149
transform 1 0 37352 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1644511149
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_41
timestamp 1644511149
transform 1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_60
timestamp 1644511149
transform 1 0 6624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_68
timestamp 1644511149
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1644511149
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_95
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1644511149
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1644511149
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1644511149
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1644511149
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_136
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_144
timestamp 1644511149
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1644511149
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1644511149
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_176
timestamp 1644511149
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_232
timestamp 1644511149
transform 1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1644511149
transform 1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1644511149
transform 1 0 24196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_259
timestamp 1644511149
transform 1 0 24932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_265
timestamp 1644511149
transform 1 0 25484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1644511149
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1644511149
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_307
timestamp 1644511149
transform 1 0 29348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_315
timestamp 1644511149
transform 1 0 30084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1644511149
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1644511149
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_344
timestamp 1644511149
transform 1 0 32752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_355
timestamp 1644511149
transform 1 0 33764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_363
timestamp 1644511149
transform 1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_370
timestamp 1644511149
transform 1 0 35144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_377
timestamp 1644511149
transform 1 0 35788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1644511149
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1644511149
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1644511149
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1644511149
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1644511149
transform 1 0 7820 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1644511149
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_119
timestamp 1644511149
transform 1 0 12052 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1644511149
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1644511149
transform 1 0 14536 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_156
timestamp 1644511149
transform 1 0 15456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1644511149
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_200
timestamp 1644511149
transform 1 0 19504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_222
timestamp 1644511149
transform 1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1644511149
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_275
timestamp 1644511149
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_326
timestamp 1644511149
transform 1 0 31096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_339
timestamp 1644511149
transform 1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_351
timestamp 1644511149
transform 1 0 33396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1644511149
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_393
timestamp 1644511149
transform 1 0 37260 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1644511149
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 1644511149
transform 1 0 4324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_64
timestamp 1644511149
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_72
timestamp 1644511149
transform 1 0 7728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1644511149
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_87
timestamp 1644511149
transform 1 0 9108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_101
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1644511149
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_150
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1644511149
transform 1 0 17296 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_199
timestamp 1644511149
transform 1 0 19412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1644511149
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_284
timestamp 1644511149
transform 1 0 27232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_288
timestamp 1644511149
transform 1 0 27600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1644511149
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_353
timestamp 1644511149
transform 1 0 33580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_365
timestamp 1644511149
transform 1 0 34684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_380
timestamp 1644511149
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_50
timestamp 1644511149
transform 1 0 5704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1644511149
transform 1 0 6440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1644511149
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_70
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1644511149
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1644511149
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_96
timestamp 1644511149
transform 1 0 9936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_101
timestamp 1644511149
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1644511149
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1644511149
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1644511149
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1644511149
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1644511149
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1644511149
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_205
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1644511149
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_261
timestamp 1644511149
transform 1 0 25116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_267
timestamp 1644511149
transform 1 0 25668 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_273
timestamp 1644511149
transform 1 0 26220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_293
timestamp 1644511149
transform 1 0 28060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1644511149
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_317
timestamp 1644511149
transform 1 0 30268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_325
timestamp 1644511149
transform 1 0 31004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1644511149
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1644511149
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_353
timestamp 1644511149
transform 1 0 33580 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_373
timestamp 1644511149
transform 1 0 35420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_381
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_393
timestamp 1644511149
transform 1 0 37260 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1644511149
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_47
timestamp 1644511149
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1644511149
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_97
timestamp 1644511149
transform 1 0 10028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1644511149
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1644511149
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_172
timestamp 1644511149
transform 1 0 16928 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_190
timestamp 1644511149
transform 1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_212
timestamp 1644511149
transform 1 0 20608 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1644511149
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_228
timestamp 1644511149
transform 1 0 22080 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_239
timestamp 1644511149
transform 1 0 23092 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_269
timestamp 1644511149
transform 1 0 25852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_285
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_297
timestamp 1644511149
transform 1 0 28428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1644511149
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_340
timestamp 1644511149
transform 1 0 32384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_348
timestamp 1644511149
transform 1 0 33120 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_356
timestamp 1644511149
transform 1 0 33856 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_370
timestamp 1644511149
transform 1 0 35144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_377
timestamp 1644511149
transform 1 0 35788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1644511149
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1644511149
transform 1 0 11868 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_125
timestamp 1644511149
transform 1 0 12604 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_131
timestamp 1644511149
transform 1 0 13156 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1644511149
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_168
timestamp 1644511149
transform 1 0 16560 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1644511149
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1644511149
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1644511149
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1644511149
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_262
timestamp 1644511149
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1644511149
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1644511149
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_294
timestamp 1644511149
transform 1 0 28152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1644511149
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1644511149
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_334
timestamp 1644511149
transform 1 0 31832 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_342
timestamp 1644511149
transform 1 0 32568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_353
timestamp 1644511149
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_47
timestamp 1644511149
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1644511149
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1644511149
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1644511149
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_143
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1644511149
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_188
timestamp 1644511149
transform 1 0 18400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_232
timestamp 1644511149
transform 1 0 22448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1644511149
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_246
timestamp 1644511149
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_252
timestamp 1644511149
transform 1 0 24288 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_269
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 1644511149
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1644511149
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_343
timestamp 1644511149
transform 1 0 32660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_363
timestamp 1644511149
transform 1 0 34500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1644511149
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1644511149
transform 1 0 7176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_70
timestamp 1644511149
transform 1 0 7544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1644511149
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1644511149
transform 1 0 9200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1644511149
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_116
timestamp 1644511149
transform 1 0 11776 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_120
timestamp 1644511149
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1644511149
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_149
timestamp 1644511149
transform 1 0 14812 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_161
timestamp 1644511149
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1644511149
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_205
timestamp 1644511149
transform 1 0 19964 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_211
timestamp 1644511149
transform 1 0 20516 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_228
timestamp 1644511149
transform 1 0 22080 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_260
timestamp 1644511149
transform 1 0 25024 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_282
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_290
timestamp 1644511149
transform 1 0 27784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1644511149
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1644511149
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_323
timestamp 1644511149
transform 1 0 30820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_343
timestamp 1644511149
transform 1 0 32660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_94
timestamp 1644511149
transform 1 0 9752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1644511149
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1644511149
transform 1 0 18032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_232
timestamp 1644511149
transform 1 0 22448 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_240
timestamp 1644511149
transform 1 0 23184 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1644511149
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1644511149
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1644511149
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_310
timestamp 1644511149
transform 1 0 29624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1644511149
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_325
timestamp 1644511149
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1644511149
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_344
timestamp 1644511149
transform 1 0 32752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_350
timestamp 1644511149
transform 1 0 33304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_358
timestamp 1644511149
transform 1 0 34040 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_370
timestamp 1644511149
transform 1 0 35144 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_382
timestamp 1644511149
transform 1 0 36248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1644511149
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_181
timestamp 1644511149
transform 1 0 17756 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1644511149
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_239
timestamp 1644511149
transform 1 0 23092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1644511149
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1644511149
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_279
timestamp 1644511149
transform 1 0 26772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_319
timestamp 1644511149
transform 1 0 30452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_330
timestamp 1644511149
transform 1 0 31464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_338
timestamp 1644511149
transform 1 0 32200 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_350
timestamp 1644511149
transform 1 0 33304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1644511149
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_234
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1644511149
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_302
timestamp 1644511149
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_323
timestamp 1644511149
transform 1 0 30820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1644511149
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_354
timestamp 1644511149
transform 1 0 33672 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_366
timestamp 1644511149
transform 1 0 34776 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_378
timestamp 1644511149
transform 1 0 35880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1644511149
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1644511149
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_260
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_279
timestamp 1644511149
transform 1 0 26772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1644511149
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_312
timestamp 1644511149
transform 1 0 29808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1644511149
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_323
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1644511149
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_335
timestamp 1644511149
transform 1 0 31924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_347
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1644511149
transform 1 0 24840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_267
timestamp 1644511149
transform 1 0 25668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1644511149
transform 1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_300
timestamp 1644511149
transform 1 0 28704 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_312
timestamp 1644511149
transform 1 0 29808 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_324
timestamp 1644511149
transform 1 0 30912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1644511149
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_342
timestamp 1644511149
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_354
timestamp 1644511149
transform 1 0 33672 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_366
timestamp 1644511149
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_378
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1644511149
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1644511149
transform 1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1644511149
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1644511149
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_256
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_276
timestamp 1644511149
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_296
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1644511149
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_324
timestamp 1644511149
transform 1 0 30912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_344
timestamp 1644511149
transform 1 0 32752 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1644511149
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_285
timestamp 1644511149
transform 1 0 27324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_340
timestamp 1644511149
transform 1 0 32384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_352
timestamp 1644511149
transform 1 0 33488 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_364
timestamp 1644511149
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_376
timestamp 1644511149
transform 1 0 35696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1644511149
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1644511149
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_294
timestamp 1644511149
transform 1 0 28152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1644511149
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1644511149
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1644511149
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1644511149
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _424_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _425_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _426_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _427_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _428_
timestamp 1644511149
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _429_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _430_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _431_
timestamp 1644511149
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _432_
timestamp 1644511149
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _433_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _434_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _435_
timestamp 1644511149
transform 1 0 15272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _436_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _437_
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _438_
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _439_
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _440_
timestamp 1644511149
transform 1 0 7912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _441_
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _442_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _443_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _444_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _445_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _446_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _447_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _448_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _449_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _450_
timestamp 1644511149
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _451_
timestamp 1644511149
transform 1 0 14168 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _452_
timestamp 1644511149
transform 1 0 13156 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _453_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _454_
timestamp 1644511149
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _455_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _456_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18768 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _457_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _458_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _459_
timestamp 1644511149
transform 1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _460_
timestamp 1644511149
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _461_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _462_
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_4  _463_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _464_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_1  _465_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _466_
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _467_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _468_
timestamp 1644511149
transform 1 0 18492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _469_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _470_
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _471_
timestamp 1644511149
transform 1 0 26312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _472_
timestamp 1644511149
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _473_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _474_
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _475_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _476_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _477_
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _478_
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _479_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _480_
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _481_
timestamp 1644511149
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _482_
timestamp 1644511149
transform 1 0 20056 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _483_
timestamp 1644511149
transform 1 0 24104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _484_
timestamp 1644511149
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _485_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _486_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _487_
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _488_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _489_
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _490_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _491_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _492_
timestamp 1644511149
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _493_
timestamp 1644511149
transform 1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp 1644511149
transform 1 0 29716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _495_
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _496_
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _497_
timestamp 1644511149
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _498_
timestamp 1644511149
transform 1 0 22448 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _499_
timestamp 1644511149
transform 1 0 23092 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp 1644511149
transform 1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _501_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _502_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _503_
timestamp 1644511149
transform 1 0 18768 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _504_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _505_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _506_
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _507_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _508_
timestamp 1644511149
transform 1 0 26680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _509_
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a221oi_2  _510_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _511_
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _512_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _513_
timestamp 1644511149
transform 1 0 23460 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _514_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _515_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _516_
timestamp 1644511149
transform 1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _517_
timestamp 1644511149
transform 1 0 24564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _518_
timestamp 1644511149
transform 1 0 28612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _519_
timestamp 1644511149
transform 1 0 25852 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _522_
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _523_
timestamp 1644511149
transform 1 0 25668 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _524_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1644511149
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _526_
timestamp 1644511149
transform 1 0 26128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _527_
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _528_
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1644511149
transform 1 0 29072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _530_
timestamp 1644511149
transform 1 0 28060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _531_
timestamp 1644511149
transform 1 0 27784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1644511149
transform 1 0 30176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _533_
timestamp 1644511149
transform 1 0 27508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _534_
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _535_
timestamp 1644511149
transform 1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _536_
timestamp 1644511149
transform 1 0 29624 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _537_
timestamp 1644511149
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _538_
timestamp 1644511149
transform 1 0 27968 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _539_
timestamp 1644511149
transform 1 0 28888 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1644511149
transform 1 0 34224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _541_
timestamp 1644511149
transform 1 0 31464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _542_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _543_
timestamp 1644511149
transform 1 0 28704 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _544_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1644511149
transform 1 0 33304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _546_
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _547_
timestamp 1644511149
transform 1 0 33948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1644511149
transform 1 0 35604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _549_
timestamp 1644511149
transform 1 0 34132 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _550_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _552_
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _553_
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp 1644511149
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _555_
timestamp 1644511149
transform 1 0 31372 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _556_
timestamp 1644511149
transform 1 0 31832 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _557_
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _559_
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _560_
timestamp 1644511149
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _561_
timestamp 1644511149
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _562_
timestamp 1644511149
transform 1 0 35144 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _563_
timestamp 1644511149
transform 1 0 35512 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1644511149
transform 1 0 36248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _566_
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _567_
timestamp 1644511149
transform 1 0 32568 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _568_
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1644511149
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _570_
timestamp 1644511149
transform 1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _571_
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _573_
timestamp 1644511149
transform 1 0 34868 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 1644511149
transform 1 0 35696 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1644511149
transform 1 0 36524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _576_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _577_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1840 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _578_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _579_
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _580_
timestamp 1644511149
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _582_
timestamp 1644511149
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _583_
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _584_
timestamp 1644511149
transform 1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _585_
timestamp 1644511149
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _586_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _587_
timestamp 1644511149
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _588_
timestamp 1644511149
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _589_
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _590_
timestamp 1644511149
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _591_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _592_
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _593_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _594_
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _595_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19320 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _596_
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _597_
timestamp 1644511149
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _598_
timestamp 1644511149
transform 1 0 18952 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _599_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _600_
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _601_
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _602_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _603_
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _604_
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _605_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _606_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _607_
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _608_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _609_
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _610_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _611_
timestamp 1644511149
transform 1 0 22724 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _612_
timestamp 1644511149
transform 1 0 28520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _613_
timestamp 1644511149
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _614_
timestamp 1644511149
transform 1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _615_
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _616_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _617_
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _618_
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _619_
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _620_
timestamp 1644511149
transform 1 0 22448 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _621_
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _622_
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _624_
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _625_
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _626_
timestamp 1644511149
transform 1 0 23000 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _627_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _628_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _630_
timestamp 1644511149
transform 1 0 12420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _631_
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _632_
timestamp 1644511149
transform 1 0 25576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _633_
timestamp 1644511149
transform 1 0 24656 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _634_
timestamp 1644511149
transform 1 0 25024 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _635_
timestamp 1644511149
transform 1 0 26312 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _636_
timestamp 1644511149
transform 1 0 25392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _637_
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _638_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _639_
timestamp 1644511149
transform 1 0 26036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _640_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _641_
timestamp 1644511149
transform 1 0 26128 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _642_
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _643_
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _644_
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _645_
timestamp 1644511149
transform 1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _646_
timestamp 1644511149
transform 1 0 27416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _647_
timestamp 1644511149
transform 1 0 26956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _648_
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _649_
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _650_
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _651_
timestamp 1644511149
transform 1 0 27232 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _652_
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _653_
timestamp 1644511149
transform 1 0 28704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _654_
timestamp 1644511149
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _655_
timestamp 1644511149
transform 1 0 28244 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _656_
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _657_
timestamp 1644511149
transform 1 0 28612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _658_
timestamp 1644511149
transform 1 0 27232 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _660_
timestamp 1644511149
transform 1 0 29900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _661_
timestamp 1644511149
transform 1 0 30544 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _662_
timestamp 1644511149
transform 1 0 30636 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _663_
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _664_
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _665_
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _666_
timestamp 1644511149
transform 1 0 30544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _667_
timestamp 1644511149
transform 1 0 30544 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _668_
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _669_
timestamp 1644511149
transform 1 0 30176 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _670_
timestamp 1644511149
transform 1 0 30820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _671_
timestamp 1644511149
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _672_
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _673_
timestamp 1644511149
transform 1 0 31004 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _674_
timestamp 1644511149
transform 1 0 30912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _675_
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _676_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _677_
timestamp 1644511149
transform 1 0 30544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _678_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _679_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _680_
timestamp 1644511149
transform 1 0 33028 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _681_
timestamp 1644511149
transform 1 0 31832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _682_
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _683_
timestamp 1644511149
transform 1 0 34224 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _684_
timestamp 1644511149
transform 1 0 32752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _685_
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _686_
timestamp 1644511149
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _687_
timestamp 1644511149
transform 1 0 33396 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _688_
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _689_
timestamp 1644511149
transform 1 0 32660 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _690_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _691_
timestamp 1644511149
transform 1 0 33120 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _692_
timestamp 1644511149
transform 1 0 32200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1644511149
transform 1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _694_
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _695_
timestamp 1644511149
transform 1 0 33764 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _696_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _697_
timestamp 1644511149
transform 1 0 31832 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _698_
timestamp 1644511149
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _699_
timestamp 1644511149
transform 1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _700_
timestamp 1644511149
transform 1 0 33948 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _701_
timestamp 1644511149
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _702_
timestamp 1644511149
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _703_
timestamp 1644511149
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _704_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _705_
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _706_
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _707_
timestamp 1644511149
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _708_
timestamp 1644511149
transform 1 0 16560 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _709_
timestamp 1644511149
transform 1 0 9476 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _710_
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _711_
timestamp 1644511149
transform 1 0 9200 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _712_
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _713_
timestamp 1644511149
transform 1 0 9568 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _714_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _715_
timestamp 1644511149
transform 1 0 11592 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _716_
timestamp 1644511149
transform 1 0 10764 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _717_
timestamp 1644511149
transform 1 0 11592 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _718_
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _719_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _720_
timestamp 1644511149
transform 1 0 9568 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _721_
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _722_
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _723_
timestamp 1644511149
transform 1 0 5152 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _724_
timestamp 1644511149
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _725_
timestamp 1644511149
transform 1 0 6532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _726_
timestamp 1644511149
transform 1 0 7728 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _727_
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _728_
timestamp 1644511149
transform 1 0 6164 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _729_
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _730_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _731_
timestamp 1644511149
transform 1 0 6716 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _732_
timestamp 1644511149
transform 1 0 6716 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _733_
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _734_
timestamp 1644511149
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _735_
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _736_
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _737_
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _738_
timestamp 1644511149
transform 1 0 7636 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _739_
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _740_
timestamp 1644511149
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _741_
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _742_
timestamp 1644511149
transform 1 0 7544 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _743_
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _744_
timestamp 1644511149
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _745_
timestamp 1644511149
transform 1 0 9108 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _746_
timestamp 1644511149
transform 1 0 9752 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _747_
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _748_
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _749_
timestamp 1644511149
transform 1 0 9384 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _750_
timestamp 1644511149
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _751_
timestamp 1644511149
transform 1 0 11316 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _752_
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _753_
timestamp 1644511149
transform 1 0 6900 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _754_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _755_
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _756_
timestamp 1644511149
transform 1 0 7912 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1644511149
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _758_
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _759_
timestamp 1644511149
transform 1 0 6992 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _761_
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp 1644511149
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp 1644511149
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _764_
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _765_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _766_
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _767_
timestamp 1644511149
transform 1 0 10212 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _768_
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _769_
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _770_
timestamp 1644511149
transform 1 0 14260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _771_
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _772_
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _773_
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _774_
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _775_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _776_
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _777_
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _778_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _779_
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _780_
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _781_
timestamp 1644511149
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _782_
timestamp 1644511149
transform 1 0 14904 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _783_
timestamp 1644511149
transform 1 0 14628 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _784_
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _785_
timestamp 1644511149
transform 1 0 12696 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _786_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _787_
timestamp 1644511149
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _788_
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _789_
timestamp 1644511149
transform 1 0 12052 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _790_
timestamp 1644511149
transform 1 0 17572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _791_
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _792_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _793_
timestamp 1644511149
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _794_
timestamp 1644511149
transform 1 0 12972 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _795_
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _796_
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _797_
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _798_
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _799_
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _800_
timestamp 1644511149
transform 1 0 13340 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _801_
timestamp 1644511149
transform 1 0 14536 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _802_
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _803_
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _804_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _805_
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _806_
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _807_
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _808_
timestamp 1644511149
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _809_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _810_
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _811_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _812_
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _813_
timestamp 1644511149
transform 1 0 14444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _814_
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _815_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _816_
timestamp 1644511149
transform 1 0 16468 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _817_
timestamp 1644511149
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _818_
timestamp 1644511149
transform 1 0 26772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _819_
timestamp 1644511149
transform 1 0 28888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _820_
timestamp 1644511149
transform 1 0 16928 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _821_
timestamp 1644511149
transform 1 0 20976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _822_
timestamp 1644511149
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _823_
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _824_
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _825_
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _826_
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _827_
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _828_
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _829_
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _830_
timestamp 1644511149
transform 1 0 20976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _831_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _832_
timestamp 1644511149
transform 1 0 21896 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _833_
timestamp 1644511149
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _834_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _835_
timestamp 1644511149
transform 1 0 22356 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _836_
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _837_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _838_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _839_
timestamp 1644511149
transform 1 0 33488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _840_
timestamp 1644511149
transform 1 0 30912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _841_
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _842_
timestamp 1644511149
transform 1 0 23368 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _843_
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _844_
timestamp 1644511149
transform 1 0 28428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _845_
timestamp 1644511149
transform 1 0 33488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _846_
timestamp 1644511149
transform 1 0 25852 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _847_
timestamp 1644511149
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _848_
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _849_
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _850_
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _851_
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _852_
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _853_
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _854_
timestamp 1644511149
transform 1 0 27600 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _855_
timestamp 1644511149
transform 1 0 35880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _856_
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _857_
timestamp 1644511149
transform 1 0 27784 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _858_
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _859_
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _860_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _861_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _862_
timestamp 1644511149
transform 1 0 35328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _863_
timestamp 1644511149
transform 1 0 36524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _864_
timestamp 1644511149
transform 1 0 33856 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _865_
timestamp 1644511149
transform 1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _866_
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _867_
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _868_
timestamp 1644511149
transform 1 0 35972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _869_
timestamp 1644511149
transform 1 0 35788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _870_
timestamp 1644511149
transform 1 0 34776 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _871_
timestamp 1644511149
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _872_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _873_
timestamp 1644511149
transform 1 0 32660 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _874_
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _875_
timestamp 1644511149
transform 1 0 28060 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _876_
timestamp 1644511149
transform 1 0 35512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _877_
timestamp 1644511149
transform 1 0 36156 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _878_
timestamp 1644511149
transform 1 0 35512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _879_
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _880_
timestamp 1644511149
transform 1 0 16744 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _881_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1644511149
transform 1 0 17940 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1644511149
transform 1 0 20608 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1644511149
transform 1 0 21620 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1644511149
transform 1 0 24196 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1644511149
transform 1 0 24380 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1644511149
transform 1 0 25576 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1644511149
transform 1 0 26864 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _900_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1644511149
transform 1 0 27508 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1644511149
transform 1 0 29532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1644511149
transform 1 0 29348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1644511149
transform 1 0 32200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1644511149
transform 1 0 30176 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1644511149
transform 1 0 31280 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1644511149
transform 1 0 31188 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1644511149
transform 1 0 33028 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1644511149
transform 1 0 34868 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1644511149
transform 1 0 32568 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1644511149
transform 1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 1644511149
transform 1 0 9108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 1644511149
transform 1 0 12328 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 1644511149
transform 1 0 4324 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 1644511149
transform 1 0 5152 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 1644511149
transform 1 0 4416 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 1644511149
transform 1 0 5244 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _923_
timestamp 1644511149
transform 1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 1644511149
transform 1 0 6624 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 1644511149
transform 1 0 7544 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1644511149
transform 1 0 6808 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1644511149
transform 1 0 9200 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1644511149
transform 1 0 10764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1644511149
transform 1 0 11316 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 1644511149
transform 1 0 12696 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 1644511149
transform 1 0 14444 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _940_
timestamp 1644511149
transform 1 0 14352 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _941_
timestamp 1644511149
transform 1 0 16376 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _942_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _943_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _944_
timestamp 1644511149
transform 1 0 15916 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _945_
timestamp 1644511149
transform 1 0 15088 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _946_
timestamp 1644511149
transform 1 0 16744 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _947_
timestamp 1644511149
transform 1 0 18400 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _948_
timestamp 1644511149
transform 1 0 22448 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 1644511149
transform 1 0 22172 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 1644511149
transform 1 0 20516 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 1644511149
transform 1 0 22264 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 1644511149
transform 1 0 23644 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _959_
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 1644511149
transform 1 0 24932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 1644511149
transform 1 0 26496 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _963_
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _964_
timestamp 1644511149
transform 1 0 27048 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _965_
timestamp 1644511149
transform 1 0 29072 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _966_
timestamp 1644511149
transform 1 0 27232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _967_
timestamp 1644511149
transform 1 0 30728 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _968_
timestamp 1644511149
transform 1 0 27600 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _969_
timestamp 1644511149
transform 1 0 29808 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _970_
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _971_
timestamp 1644511149
transform 1 0 29624 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _972_
timestamp 1644511149
transform 1 0 31648 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _973_
timestamp 1644511149
transform 1 0 29808 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _974_
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _975_
timestamp 1644511149
transform 1 0 32384 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _976_
timestamp 1644511149
transform 1 0 32200 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _977_
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _978_
timestamp 1644511149
transform 1 0 34684 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _979_
timestamp 1644511149
transform 1 0 19228 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _980_
timestamp 1644511149
transform 1 0 16836 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _981__69 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _982__70
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_CLK
timestamp 1644511149
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_CLK
timestamp 1644511149
transform 1 0 28796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_CLK
timestamp 1644511149
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_CLK
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_CLK
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_CLK
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_CLK
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_CLK
timestamp 1644511149
transform 1 0 15824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_CLK
timestamp 1644511149
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_CLK
timestamp 1644511149
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_CLK
timestamp 1644511149
transform 1 0 30636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_CLK
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_CLK
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_CLK
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1644511149
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1644511149
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1644511149
transform 1 0 35696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1644511149
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1644511149
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 25484 0 -1 6528
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 570 0 626 800 6 RST_N
port 1 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 slave_ack_o
port 2 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 slave_adr_i[0]
port 3 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 slave_adr_i[10]
port 4 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 slave_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 slave_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 slave_adr_i[13]
port 7 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 slave_adr_i[14]
port 8 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 slave_adr_i[15]
port 9 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 slave_adr_i[16]
port 10 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 slave_adr_i[17]
port 11 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 slave_adr_i[18]
port 12 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 slave_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 slave_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 slave_adr_i[20]
port 15 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 slave_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 slave_adr_i[22]
port 17 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 slave_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 slave_adr_i[24]
port 19 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 slave_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 slave_adr_i[26]
port 21 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 slave_adr_i[27]
port 22 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 slave_adr_i[28]
port 23 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 slave_adr_i[29]
port 24 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 slave_adr_i[2]
port 25 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 slave_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 slave_adr_i[31]
port 27 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 slave_adr_i[3]
port 28 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 slave_adr_i[4]
port 29 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 slave_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 slave_adr_i[6]
port 31 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 slave_adr_i[7]
port 32 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 slave_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 slave_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 938 0 994 800 6 slave_cyc_i
port 35 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 slave_dat_i[0]
port 36 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 slave_dat_i[10]
port 37 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 slave_dat_i[11]
port 38 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 slave_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 slave_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 slave_dat_i[14]
port 41 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 slave_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 slave_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 slave_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 slave_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 slave_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 slave_dat_i[1]
port 47 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 slave_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 slave_dat_i[21]
port 49 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 slave_dat_i[22]
port 50 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 slave_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 slave_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 slave_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 slave_dat_i[26]
port 54 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 slave_dat_i[27]
port 55 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 slave_dat_i[28]
port 56 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 slave_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 slave_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 slave_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 slave_dat_i[31]
port 60 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 slave_dat_i[3]
port 61 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 slave_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 slave_dat_i[5]
port 63 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 slave_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 slave_dat_i[7]
port 65 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 slave_dat_i[8]
port 66 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 slave_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 slave_dat_o[0]
port 68 nsew signal tristate
rlabel metal2 s 24122 0 24178 800 6 slave_dat_o[10]
port 69 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 slave_dat_o[11]
port 70 nsew signal tristate
rlabel metal2 s 25594 0 25650 800 6 slave_dat_o[12]
port 71 nsew signal tristate
rlabel metal2 s 26330 0 26386 800 6 slave_dat_o[13]
port 72 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 slave_dat_o[14]
port 73 nsew signal tristate
rlabel metal2 s 27802 0 27858 800 6 slave_dat_o[15]
port 74 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 slave_dat_o[16]
port 75 nsew signal tristate
rlabel metal2 s 29366 0 29422 800 6 slave_dat_o[17]
port 76 nsew signal tristate
rlabel metal2 s 30102 0 30158 800 6 slave_dat_o[18]
port 77 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 slave_dat_o[19]
port 78 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 slave_dat_o[1]
port 79 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 slave_dat_o[20]
port 80 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 slave_dat_o[21]
port 81 nsew signal tristate
rlabel metal2 s 33046 0 33102 800 6 slave_dat_o[22]
port 82 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 slave_dat_o[23]
port 83 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 slave_dat_o[24]
port 84 nsew signal tristate
rlabel metal2 s 35346 0 35402 800 6 slave_dat_o[25]
port 85 nsew signal tristate
rlabel metal2 s 36082 0 36138 800 6 slave_dat_o[26]
port 86 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 slave_dat_o[27]
port 87 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 slave_dat_o[28]
port 88 nsew signal tristate
rlabel metal2 s 38290 0 38346 800 6 slave_dat_o[29]
port 89 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 slave_dat_o[2]
port 90 nsew signal tristate
rlabel metal2 s 39026 0 39082 800 6 slave_dat_o[30]
port 91 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 slave_dat_o[31]
port 92 nsew signal tristate
rlabel metal2 s 18878 0 18934 800 6 slave_dat_o[3]
port 93 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 slave_dat_o[4]
port 94 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 slave_dat_o[5]
port 95 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 slave_dat_o[6]
port 96 nsew signal tristate
rlabel metal2 s 21822 0 21878 800 6 slave_dat_o[7]
port 97 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 slave_dat_o[8]
port 98 nsew signal tristate
rlabel metal2 s 23386 0 23442 800 6 slave_dat_o[9]
port 99 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 slave_err_o
port 100 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 slave_rty_o
port 101 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 slave_sel_i[0]
port 102 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 slave_sel_i[1]
port 103 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 slave_sel_i[2]
port 104 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 slave_sel_i[3]
port 105 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 slave_stb_i
port 106 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 slave_we_i
port 107 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 108 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 108 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 109 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
