magic
tech sky130A
magscale 1 2
timestamp 1647707505
<< viali >>
rect 15209 47209 15243 47243
rect 25237 47209 25271 47243
rect 35265 47209 35299 47243
rect 5089 47005 5123 47039
rect 15025 47005 15059 47039
rect 25053 47005 25087 47039
rect 35081 47005 35115 47039
rect 5273 46869 5307 46903
rect 19809 46665 19843 46699
rect 19993 46529 20027 46563
rect 19441 30685 19475 30719
rect 19257 30549 19291 30583
rect 19248 30277 19282 30311
rect 17141 30209 17175 30243
rect 17408 30209 17442 30243
rect 18981 30209 19015 30243
rect 18521 30005 18555 30039
rect 20361 30005 20395 30039
rect 18429 29801 18463 29835
rect 21005 29801 21039 29835
rect 15761 29665 15795 29699
rect 19809 29665 19843 29699
rect 20637 29665 20671 29699
rect 17601 29597 17635 29631
rect 17785 29597 17819 29631
rect 17969 29597 18003 29631
rect 18613 29597 18647 29631
rect 19993 29597 20027 29631
rect 20821 29597 20855 29631
rect 16028 29529 16062 29563
rect 17141 29461 17175 29495
rect 20177 29461 20211 29495
rect 16681 29257 16715 29291
rect 18429 29257 18463 29291
rect 19441 29257 19475 29291
rect 21833 29257 21867 29291
rect 19165 29189 19199 29223
rect 20168 29189 20202 29223
rect 15945 29121 15979 29155
rect 16865 29121 16899 29155
rect 17877 29121 17911 29155
rect 18061 29121 18095 29155
rect 18153 29121 18187 29155
rect 18291 29121 18325 29155
rect 18889 29121 18923 29155
rect 19073 29121 19107 29155
rect 19257 29121 19291 29155
rect 22017 29121 22051 29155
rect 19901 29053 19935 29087
rect 21281 28985 21315 29019
rect 15761 28917 15795 28951
rect 19809 28713 19843 28747
rect 22661 28713 22695 28747
rect 15853 28577 15887 28611
rect 22293 28577 22327 28611
rect 16120 28509 16154 28543
rect 17693 28509 17727 28543
rect 18061 28509 18095 28543
rect 19257 28509 19291 28543
rect 19625 28509 19659 28543
rect 20453 28509 20487 28543
rect 22477 28509 22511 28543
rect 17877 28441 17911 28475
rect 17969 28441 18003 28475
rect 19441 28441 19475 28475
rect 19533 28441 19567 28475
rect 20720 28441 20754 28475
rect 17233 28373 17267 28407
rect 18245 28373 18279 28407
rect 21833 28373 21867 28407
rect 15853 28169 15887 28203
rect 17049 28169 17083 28203
rect 17693 28169 17727 28203
rect 18889 28169 18923 28203
rect 20637 28169 20671 28203
rect 21097 28169 21131 28203
rect 15025 28033 15059 28067
rect 15669 28033 15703 28067
rect 16865 28033 16899 28067
rect 18061 28033 18095 28067
rect 19257 28033 19291 28067
rect 20085 28033 20119 28067
rect 20269 28033 20303 28067
rect 20361 28033 20395 28067
rect 20453 28033 20487 28067
rect 21281 28033 21315 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22661 28033 22695 28067
rect 22928 28033 22962 28067
rect 24768 28033 24802 28067
rect 15485 27965 15519 27999
rect 16681 27965 16715 27999
rect 18153 27965 18187 27999
rect 18337 27965 18371 27999
rect 19349 27965 19383 27999
rect 19533 27965 19567 27999
rect 24501 27965 24535 27999
rect 14841 27897 14875 27931
rect 21833 27829 21867 27863
rect 24041 27829 24075 27863
rect 25881 27829 25915 27863
rect 20453 27625 20487 27659
rect 17233 27557 17267 27591
rect 19257 27557 19291 27591
rect 24409 27557 24443 27591
rect 15945 27489 15979 27523
rect 17877 27489 17911 27523
rect 19809 27489 19843 27523
rect 21097 27489 21131 27523
rect 22109 27489 22143 27523
rect 14105 27421 14139 27455
rect 16221 27421 16255 27455
rect 17417 27421 17451 27455
rect 18153 27421 18187 27455
rect 19717 27421 19751 27455
rect 20913 27421 20947 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 14350 27353 14384 27387
rect 22376 27353 22410 27387
rect 15485 27285 15519 27319
rect 19625 27285 19659 27319
rect 20821 27285 20855 27319
rect 23489 27285 23523 27319
rect 25329 27285 25363 27319
rect 13369 27081 13403 27115
rect 17233 27081 17267 27115
rect 19257 27081 19291 27115
rect 20545 27081 20579 27115
rect 16957 27013 16991 27047
rect 19717 27013 19751 27047
rect 25513 27013 25547 27047
rect 13553 26945 13587 26979
rect 14197 26945 14231 26979
rect 14657 26945 14691 26979
rect 14913 26945 14947 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 17049 26945 17083 26979
rect 18245 26945 18279 26979
rect 19625 26945 19659 26979
rect 20453 26945 20487 26979
rect 20637 26945 20671 26979
rect 21097 26945 21131 26979
rect 21281 26945 21315 26979
rect 22109 26945 22143 26979
rect 22569 26945 22603 26979
rect 23949 26945 23983 26979
rect 24409 26945 24443 26979
rect 25329 26945 25363 26979
rect 25605 26945 25639 26979
rect 26065 26945 26099 26979
rect 27241 26945 27275 26979
rect 17969 26877 18003 26911
rect 19901 26877 19935 26911
rect 21189 26877 21223 26911
rect 22845 26877 22879 26911
rect 24133 26877 24167 26911
rect 24225 26877 24259 26911
rect 26985 26877 27019 26911
rect 14013 26809 14047 26843
rect 24041 26809 24075 26843
rect 26249 26809 26283 26843
rect 16037 26741 16071 26775
rect 23765 26741 23799 26775
rect 25145 26741 25179 26775
rect 28365 26741 28399 26775
rect 15669 26537 15703 26571
rect 16497 26537 16531 26571
rect 17049 26537 17083 26571
rect 18521 26537 18555 26571
rect 19349 26537 19383 26571
rect 21281 26537 21315 26571
rect 22201 26537 22235 26571
rect 23673 26537 23707 26571
rect 23857 26537 23891 26571
rect 24409 26537 24443 26571
rect 25145 26537 25179 26571
rect 26893 26537 26927 26571
rect 14841 26469 14875 26503
rect 25513 26469 25547 26503
rect 17693 26401 17727 26435
rect 21005 26401 21039 26435
rect 22017 26401 22051 26435
rect 25421 26401 25455 26435
rect 28181 26401 28215 26435
rect 12817 26333 12851 26367
rect 13001 26333 13035 26367
rect 14289 26333 14323 26367
rect 14657 26333 14691 26367
rect 15393 26333 15427 26367
rect 15485 26333 15519 26367
rect 16129 26333 16163 26367
rect 16313 26333 16347 26367
rect 18521 26333 18555 26367
rect 18705 26333 18739 26367
rect 19349 26333 19383 26367
rect 19533 26333 19567 26367
rect 20085 26333 20119 26367
rect 20269 26333 20303 26367
rect 20913 26333 20947 26367
rect 21925 26333 21959 26367
rect 22753 26333 22787 26367
rect 24685 26333 24719 26367
rect 25329 26333 25363 26367
rect 25605 26333 25639 26367
rect 25789 26333 25823 26367
rect 26249 26333 26283 26367
rect 26433 26333 26467 26367
rect 27077 26333 27111 26367
rect 27169 26333 27203 26367
rect 27353 26333 27387 26367
rect 27445 26333 27479 26367
rect 27906 26333 27940 26367
rect 27997 26333 28031 26367
rect 14473 26265 14507 26299
rect 14565 26265 14599 26299
rect 17417 26265 17451 26299
rect 17509 26265 17543 26299
rect 23489 26265 23523 26299
rect 23705 26265 23739 26299
rect 24409 26265 24443 26299
rect 26341 26265 26375 26299
rect 13185 26197 13219 26231
rect 20269 26197 20303 26231
rect 22937 26197 22971 26231
rect 24593 26197 24627 26231
rect 28181 26197 28215 26231
rect 14105 25993 14139 26027
rect 21005 25993 21039 26027
rect 27353 25993 27387 26027
rect 14565 25925 14599 25959
rect 24593 25925 24627 25959
rect 26433 25925 26467 25959
rect 27813 25925 27847 25959
rect 27997 25925 28031 25959
rect 12429 25857 12463 25891
rect 14473 25857 14507 25891
rect 16865 25857 16899 25891
rect 17049 25857 17083 25891
rect 17693 25857 17727 25891
rect 18429 25857 18463 25891
rect 18613 25857 18647 25891
rect 19257 25857 19291 25891
rect 19441 25857 19475 25891
rect 19901 25857 19935 25891
rect 20085 25857 20119 25891
rect 20637 25857 20671 25891
rect 20821 25857 20855 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22661 25857 22695 25891
rect 22845 25857 22879 25891
rect 23673 25857 23707 25891
rect 24317 25857 24351 25891
rect 24409 25857 24443 25891
rect 25329 25857 25363 25891
rect 25421 25857 25455 25891
rect 25513 25857 25547 25891
rect 25697 25857 25731 25891
rect 26249 25857 26283 25891
rect 27169 25857 27203 25891
rect 28089 25857 28123 25891
rect 28549 25857 28583 25891
rect 28733 25857 28767 25891
rect 31125 25857 31159 25891
rect 31309 25857 31343 25891
rect 12173 25789 12207 25823
rect 14749 25789 14783 25823
rect 15301 25789 15335 25823
rect 15577 25789 15611 25823
rect 16681 25789 16715 25823
rect 24593 25789 24627 25823
rect 26985 25789 27019 25823
rect 19257 25721 19291 25755
rect 27813 25721 27847 25755
rect 13553 25653 13587 25687
rect 17509 25653 17543 25687
rect 18429 25653 18463 25687
rect 19901 25653 19935 25687
rect 20821 25653 20855 25687
rect 21925 25653 21959 25687
rect 25053 25653 25087 25687
rect 28549 25653 28583 25687
rect 31217 25653 31251 25687
rect 12173 25449 12207 25483
rect 20545 25449 20579 25483
rect 23857 25449 23891 25483
rect 25053 25449 25087 25483
rect 19257 25381 19291 25415
rect 20729 25381 20763 25415
rect 13461 25313 13495 25347
rect 16313 25313 16347 25347
rect 20453 25313 20487 25347
rect 21189 25313 21223 25347
rect 22569 25313 22603 25347
rect 23029 25313 23063 25347
rect 25605 25313 25639 25347
rect 12357 25245 12391 25279
rect 14657 25245 14691 25279
rect 14933 25245 14967 25279
rect 16580 25245 16614 25279
rect 18245 25245 18279 25279
rect 18429 25245 18463 25279
rect 19257 25245 19291 25279
rect 19435 25245 19469 25279
rect 20361 25245 20395 25279
rect 21465 25245 21499 25279
rect 22661 25245 22695 25279
rect 23489 25245 23523 25279
rect 24961 25245 24995 25279
rect 25145 25245 25179 25279
rect 25861 25245 25895 25279
rect 27629 25245 27663 25279
rect 27896 25245 27930 25279
rect 29837 25245 29871 25279
rect 31677 25245 31711 25279
rect 13277 25177 13311 25211
rect 23673 25177 23707 25211
rect 30104 25177 30138 25211
rect 31922 25177 31956 25211
rect 12817 25109 12851 25143
rect 13185 25109 13219 25143
rect 17693 25109 17727 25143
rect 18337 25109 18371 25143
rect 26985 25109 27019 25143
rect 29009 25109 29043 25143
rect 31217 25109 31251 25143
rect 33057 25109 33091 25143
rect 17325 24905 17359 24939
rect 18705 24905 18739 24939
rect 22063 24905 22097 24939
rect 26265 24905 26299 24939
rect 27813 24905 27847 24939
rect 28457 24905 28491 24939
rect 13277 24837 13311 24871
rect 14473 24837 14507 24871
rect 26065 24837 26099 24871
rect 13093 24769 13127 24803
rect 13369 24769 13403 24803
rect 13461 24769 13495 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 18521 24769 18555 24803
rect 19625 24769 19659 24803
rect 20637 24769 20671 24803
rect 20821 24769 20855 24803
rect 21833 24769 21867 24803
rect 23121 24769 23155 24803
rect 24225 24769 24259 24803
rect 25237 24769 25271 24803
rect 25421 24769 25455 24803
rect 26985 24769 27019 24803
rect 27629 24769 27663 24803
rect 27905 24769 27939 24803
rect 28365 24769 28399 24803
rect 28549 24769 28583 24803
rect 29101 24769 29135 24803
rect 29368 24769 29402 24803
rect 31033 24769 31067 24803
rect 32597 24769 32631 24803
rect 32781 24769 32815 24803
rect 14565 24701 14599 24735
rect 14749 24701 14783 24735
rect 15301 24701 15335 24735
rect 15577 24701 15611 24735
rect 17417 24701 17451 24735
rect 17601 24701 17635 24735
rect 19349 24701 19383 24735
rect 23213 24701 23247 24735
rect 13645 24633 13679 24667
rect 14105 24633 14139 24667
rect 25237 24633 25271 24667
rect 26433 24633 26467 24667
rect 31217 24633 31251 24667
rect 16957 24565 16991 24599
rect 20637 24565 20671 24599
rect 21005 24565 21039 24599
rect 23121 24565 23155 24599
rect 23489 24565 23523 24599
rect 24041 24565 24075 24599
rect 26249 24565 26283 24599
rect 27077 24565 27111 24599
rect 27629 24565 27663 24599
rect 30481 24565 30515 24599
rect 32597 24565 32631 24599
rect 17877 24361 17911 24395
rect 20729 24361 20763 24395
rect 24869 24361 24903 24395
rect 25605 24361 25639 24395
rect 26341 24361 26375 24395
rect 30021 24361 30055 24395
rect 33517 24361 33551 24395
rect 19257 24293 19291 24327
rect 20913 24293 20947 24327
rect 30205 24293 30239 24327
rect 15025 24225 15059 24259
rect 21741 24225 21775 24259
rect 23673 24225 23707 24259
rect 24501 24225 24535 24259
rect 30665 24225 30699 24259
rect 12541 24157 12575 24191
rect 13001 24157 13035 24191
rect 13369 24157 13403 24191
rect 14749 24157 14783 24191
rect 16037 24157 16071 24191
rect 16313 24157 16347 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 19257 24157 19291 24191
rect 19441 24157 19475 24191
rect 19901 24157 19935 24191
rect 20085 24157 20119 24191
rect 20550 24157 20584 24191
rect 20729 24157 20763 24191
rect 22017 24157 22051 24191
rect 23489 24157 23523 24191
rect 24593 24157 24627 24191
rect 26249 24157 26283 24191
rect 27445 24157 27479 24191
rect 27712 24157 27746 24191
rect 29837 24157 29871 24191
rect 30021 24157 30055 24191
rect 30941 24157 30975 24191
rect 32137 24157 32171 24191
rect 13185 24089 13219 24123
rect 13277 24089 13311 24123
rect 17601 24089 17635 24123
rect 23581 24089 23615 24123
rect 25421 24089 25455 24123
rect 32404 24089 32438 24123
rect 12357 24021 12391 24055
rect 13553 24021 13587 24055
rect 18337 24021 18371 24055
rect 19993 24021 20027 24055
rect 23121 24021 23155 24055
rect 25621 24021 25655 24055
rect 25789 24021 25823 24055
rect 28825 24021 28859 24055
rect 13921 23817 13955 23851
rect 14289 23817 14323 23851
rect 17049 23817 17083 23851
rect 21281 23817 21315 23851
rect 22033 23817 22067 23851
rect 26985 23817 27019 23851
rect 28089 23817 28123 23851
rect 33333 23817 33367 23851
rect 12072 23749 12106 23783
rect 20453 23749 20487 23783
rect 21833 23749 21867 23783
rect 27353 23749 27387 23783
rect 29009 23749 29043 23783
rect 32873 23749 32907 23783
rect 11805 23681 11839 23715
rect 15301 23681 15335 23715
rect 17877 23681 17911 23715
rect 18061 23681 18095 23715
rect 18153 23681 18187 23715
rect 18291 23681 18325 23715
rect 19441 23681 19475 23715
rect 20269 23681 20303 23715
rect 20913 23681 20947 23715
rect 21097 23681 21131 23715
rect 22661 23681 22695 23715
rect 22845 23681 22879 23715
rect 23673 23681 23707 23715
rect 24317 23681 24351 23715
rect 25237 23681 25271 23715
rect 25421 23681 25455 23715
rect 25973 23681 26007 23715
rect 26157 23681 26191 23715
rect 27169 23681 27203 23715
rect 27445 23681 27479 23715
rect 28086 23681 28120 23715
rect 29193 23681 29227 23715
rect 29285 23681 29319 23715
rect 30297 23681 30331 23715
rect 32137 23681 32171 23715
rect 32321 23681 32355 23715
rect 32413 23681 32447 23715
rect 32689 23681 32723 23715
rect 33609 23681 33643 23715
rect 33701 23681 33735 23715
rect 33793 23681 33827 23715
rect 33953 23681 33987 23715
rect 34437 23681 34471 23715
rect 34621 23681 34655 23715
rect 14381 23613 14415 23647
rect 14565 23613 14599 23647
rect 15577 23613 15611 23647
rect 17141 23613 17175 23647
rect 17325 23613 17359 23647
rect 20085 23613 20119 23647
rect 22753 23613 22787 23647
rect 25145 23613 25179 23647
rect 25329 23613 25363 23647
rect 28549 23613 28583 23647
rect 30573 23613 30607 23647
rect 32505 23613 32539 23647
rect 13185 23545 13219 23579
rect 22201 23545 22235 23579
rect 23857 23545 23891 23579
rect 28457 23545 28491 23579
rect 16681 23477 16715 23511
rect 18429 23477 18463 23511
rect 19533 23477 19567 23511
rect 21097 23477 21131 23511
rect 22017 23477 22051 23511
rect 24409 23477 24443 23511
rect 24961 23477 24995 23511
rect 25973 23477 26007 23511
rect 27905 23477 27939 23511
rect 29009 23477 29043 23511
rect 34529 23477 34563 23511
rect 12541 23273 12575 23307
rect 17693 23273 17727 23307
rect 20453 23273 20487 23307
rect 22937 23273 22971 23307
rect 26341 23273 26375 23307
rect 30665 23273 30699 23307
rect 34805 23273 34839 23307
rect 13553 23205 13587 23239
rect 27537 23205 27571 23239
rect 31125 23205 31159 23239
rect 12173 23137 12207 23171
rect 16957 23137 16991 23171
rect 17141 23137 17175 23171
rect 18337 23137 18371 23171
rect 20453 23137 20487 23171
rect 21925 23137 21959 23171
rect 23857 23137 23891 23171
rect 30205 23137 30239 23171
rect 32505 23137 32539 23171
rect 33609 23137 33643 23171
rect 11437 23069 11471 23103
rect 11529 23069 11563 23103
rect 12357 23069 12391 23103
rect 13001 23069 13035 23103
rect 13185 23069 13219 23103
rect 13369 23069 13403 23103
rect 14657 23069 14691 23103
rect 14933 23069 14967 23103
rect 19257 23069 19291 23103
rect 19533 23069 19567 23103
rect 19625 23069 19659 23103
rect 20361 23069 20395 23103
rect 20637 23069 20671 23103
rect 21649 23069 21683 23103
rect 22937 23069 22971 23103
rect 23121 23069 23155 23103
rect 24961 23069 24995 23103
rect 25217 23069 25251 23103
rect 29929 23069 29963 23103
rect 30113 23069 30147 23103
rect 30297 23069 30331 23103
rect 30481 23069 30515 23103
rect 31401 23069 31435 23103
rect 32137 23069 32171 23103
rect 32321 23069 32355 23103
rect 32413 23069 32447 23103
rect 32689 23069 32723 23103
rect 33333 23069 33367 23103
rect 34713 23069 34747 23103
rect 13277 23001 13311 23035
rect 18061 23001 18095 23035
rect 23673 23001 23707 23035
rect 27169 23001 27203 23035
rect 28457 23001 28491 23035
rect 28641 23001 28675 23035
rect 31125 23001 31159 23035
rect 11713 22933 11747 22967
rect 16497 22933 16531 22967
rect 16865 22933 16899 22967
rect 18153 22933 18187 22967
rect 20821 22933 20855 22967
rect 27629 22933 27663 22967
rect 28825 22933 28859 22967
rect 31309 22933 31343 22967
rect 32873 22933 32907 22967
rect 14841 22729 14875 22763
rect 21189 22729 21223 22763
rect 22585 22729 22619 22763
rect 22753 22729 22787 22763
rect 25053 22729 25087 22763
rect 28825 22729 28859 22763
rect 29745 22729 29779 22763
rect 30665 22729 30699 22763
rect 32229 22729 32263 22763
rect 17500 22661 17534 22695
rect 22385 22661 22419 22695
rect 27537 22661 27571 22695
rect 30113 22661 30147 22695
rect 32597 22661 32631 22695
rect 33578 22661 33612 22695
rect 11989 22593 12023 22627
rect 12256 22593 12290 22627
rect 14013 22593 14047 22627
rect 15761 22593 15795 22627
rect 15853 22593 15887 22627
rect 17233 22593 17267 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 20177 22593 20211 22627
rect 20453 22593 20487 22627
rect 21097 22593 21131 22627
rect 21281 22593 21315 22627
rect 23305 22593 23339 22627
rect 24041 22593 24075 22627
rect 24225 22593 24259 22627
rect 24961 22593 24995 22627
rect 25605 22593 25639 22627
rect 27721 22593 27755 22627
rect 27997 22593 28031 22627
rect 28549 22593 28583 22627
rect 28733 22593 28767 22627
rect 29929 22593 29963 22627
rect 30205 22593 30239 22627
rect 30895 22593 30929 22627
rect 31030 22593 31064 22627
rect 31125 22593 31159 22627
rect 31309 22593 31343 22627
rect 32413 22593 32447 22627
rect 32689 22593 32723 22627
rect 33333 22593 33367 22627
rect 14933 22525 14967 22559
rect 15117 22525 15151 22559
rect 20361 22525 20395 22559
rect 25881 22525 25915 22559
rect 13829 22457 13863 22491
rect 19717 22457 19751 22491
rect 20637 22457 20671 22491
rect 27813 22457 27847 22491
rect 27905 22457 27939 22491
rect 13369 22389 13403 22423
rect 14473 22389 14507 22423
rect 16037 22389 16071 22423
rect 18613 22389 18647 22423
rect 19441 22389 19475 22423
rect 20453 22389 20487 22423
rect 22569 22389 22603 22423
rect 23397 22389 23431 22423
rect 24133 22389 24167 22423
rect 34713 22389 34747 22423
rect 17601 22185 17635 22219
rect 19901 22185 19935 22219
rect 25697 22185 25731 22219
rect 27813 22185 27847 22219
rect 28825 22185 28859 22219
rect 29653 22185 29687 22219
rect 30297 22185 30331 22219
rect 33609 22185 33643 22219
rect 13553 22117 13587 22151
rect 16497 22049 16531 22083
rect 18429 22049 18463 22083
rect 20913 22049 20947 22083
rect 25145 22049 25179 22083
rect 25303 22049 25337 22083
rect 25513 22049 25547 22083
rect 29837 22049 29871 22083
rect 31217 22049 31251 22083
rect 32689 22049 32723 22083
rect 32781 22049 32815 22083
rect 33793 22049 33827 22083
rect 12265 21981 12299 22015
rect 12357 21981 12391 22015
rect 13001 21981 13035 22015
rect 13185 21981 13219 22015
rect 13369 21981 13403 22015
rect 14841 21981 14875 22015
rect 15209 21981 15243 22015
rect 16221 21981 16255 22015
rect 17049 21981 17083 22015
rect 17233 21981 17267 22015
rect 17417 21981 17451 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 20177 21981 20211 22015
rect 20637 21981 20671 22015
rect 22109 21981 22143 22015
rect 24685 21981 24719 22015
rect 26433 21981 26467 22015
rect 26709 21981 26743 22015
rect 27353 21981 27387 22015
rect 27721 21981 27755 22015
rect 27997 21981 28031 22015
rect 28457 21981 28491 22015
rect 29561 21981 29595 22015
rect 30297 21981 30331 22015
rect 30481 21981 30515 22015
rect 30941 21981 30975 22015
rect 32413 21981 32447 22015
rect 32597 21981 32631 22015
rect 32965 21981 32999 22015
rect 33885 21981 33919 22015
rect 13277 21913 13311 21947
rect 15025 21913 15059 21947
rect 15117 21913 15151 21947
rect 17325 21913 17359 21947
rect 19717 21913 19751 21947
rect 22376 21913 22410 21947
rect 24501 21913 24535 21947
rect 26157 21913 26191 21947
rect 28641 21913 28675 21947
rect 29837 21913 29871 21947
rect 33609 21913 33643 21947
rect 12541 21845 12575 21879
rect 15393 21845 15427 21879
rect 15853 21845 15887 21879
rect 16313 21845 16347 21879
rect 19901 21845 19935 21879
rect 23489 21845 23523 21879
rect 26341 21845 26375 21879
rect 26525 21845 26559 21879
rect 27537 21845 27571 21879
rect 33149 21845 33183 21879
rect 34069 21845 34103 21879
rect 17141 21641 17175 21675
rect 22201 21641 22235 21675
rect 22937 21641 22971 21675
rect 24685 21641 24719 21675
rect 31217 21641 31251 21675
rect 32137 21641 32171 21675
rect 34897 21641 34931 21675
rect 21833 21573 21867 21607
rect 22033 21573 22067 21607
rect 23305 21573 23339 21607
rect 25605 21573 25639 21607
rect 26157 21573 26191 21607
rect 27169 21573 27203 21607
rect 30481 21573 30515 21607
rect 30941 21573 30975 21607
rect 31125 21573 31159 21607
rect 33762 21573 33796 21607
rect 35633 21573 35667 21607
rect 12817 21505 12851 21539
rect 13084 21505 13118 21539
rect 15005 21505 15039 21539
rect 16773 21505 16807 21539
rect 16957 21505 16991 21539
rect 18317 21505 18351 21539
rect 20453 21505 20487 21539
rect 20729 21505 20763 21539
rect 22845 21505 22879 21539
rect 23765 21505 23799 21539
rect 24593 21505 24627 21539
rect 25421 21505 25455 21539
rect 28089 21505 28123 21539
rect 28181 21505 28215 21539
rect 28273 21505 28307 21539
rect 28457 21505 28491 21539
rect 29193 21505 29227 21539
rect 29285 21505 29319 21539
rect 29377 21505 29411 21539
rect 29561 21505 29595 21539
rect 30205 21505 30239 21539
rect 31217 21505 31251 21539
rect 32321 21505 32355 21539
rect 32505 21505 32539 21539
rect 32597 21505 32631 21539
rect 35357 21505 35391 21539
rect 14749 21437 14783 21471
rect 18061 21437 18095 21471
rect 23213 21437 23247 21471
rect 25237 21437 25271 21471
rect 30481 21437 30515 21471
rect 33517 21437 33551 21471
rect 35633 21437 35667 21471
rect 23121 21369 23155 21403
rect 26341 21369 26375 21403
rect 27353 21369 27387 21403
rect 14197 21301 14231 21335
rect 16129 21301 16163 21335
rect 19441 21301 19475 21335
rect 22017 21301 22051 21335
rect 23765 21301 23799 21335
rect 27813 21301 27847 21335
rect 28917 21301 28951 21335
rect 30297 21301 30331 21335
rect 35449 21301 35483 21335
rect 13277 21097 13311 21131
rect 14749 21097 14783 21131
rect 15577 21097 15611 21131
rect 19257 21097 19291 21131
rect 20085 21097 20119 21131
rect 24777 21097 24811 21131
rect 26801 21097 26835 21131
rect 28365 21097 28399 21131
rect 29561 21097 29595 21131
rect 30665 21097 30699 21131
rect 31677 21097 31711 21131
rect 32321 21097 32355 21131
rect 33977 21097 34011 21131
rect 22661 21029 22695 21063
rect 23489 21029 23523 21063
rect 27629 21029 27663 21063
rect 31033 21029 31067 21063
rect 32689 21029 32723 21063
rect 20637 20961 20671 20995
rect 27813 20961 27847 20995
rect 29837 20961 29871 20995
rect 30757 20961 30791 20995
rect 31861 20961 31895 20995
rect 32413 20961 32447 20995
rect 33333 20961 33367 20995
rect 13461 20893 13495 20927
rect 14933 20893 14967 20927
rect 15485 20893 15519 20927
rect 16589 20893 16623 20927
rect 16773 20893 16807 20927
rect 16865 20893 16899 20927
rect 16957 20893 16991 20927
rect 17141 20893 17175 20927
rect 17325 20893 17359 20927
rect 18245 20893 18279 20927
rect 18429 20893 18463 20927
rect 18521 20893 18555 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 21741 20893 21775 20927
rect 21925 20893 21959 20927
rect 22477 20893 22511 20927
rect 23305 20893 23339 20927
rect 23581 20893 23615 20927
rect 25421 20893 25455 20927
rect 27537 20893 27571 20927
rect 28549 20893 28583 20927
rect 28643 20893 28677 20927
rect 28871 20893 28905 20927
rect 29009 20893 29043 20927
rect 29745 20893 29779 20927
rect 30205 20893 30239 20927
rect 30665 20893 30699 20927
rect 31585 20893 31619 20927
rect 32321 20893 32355 20927
rect 33149 20893 33183 20927
rect 33517 20893 33551 20927
rect 33977 20893 34011 20927
rect 34161 20893 34195 20927
rect 20453 20825 20487 20859
rect 24593 20825 24627 20859
rect 24809 20825 24843 20859
rect 25688 20825 25722 20859
rect 27813 20825 27847 20859
rect 28733 20825 28767 20859
rect 31861 20825 31895 20859
rect 18061 20757 18095 20791
rect 20545 20757 20579 20791
rect 21833 20757 21867 20791
rect 23121 20757 23155 20791
rect 24961 20757 24995 20791
rect 29929 20757 29963 20791
rect 30113 20757 30147 20791
rect 33241 20757 33275 20791
rect 33425 20757 33459 20791
rect 12909 20553 12943 20587
rect 15025 20553 15059 20587
rect 19993 20553 20027 20587
rect 26249 20553 26283 20587
rect 28457 20553 28491 20587
rect 28917 20553 28951 20587
rect 32321 20553 32355 20587
rect 32689 20553 32723 20587
rect 34897 20553 34931 20587
rect 15945 20485 15979 20519
rect 18214 20485 18248 20519
rect 20913 20485 20947 20519
rect 22017 20485 22051 20519
rect 33762 20485 33796 20519
rect 12817 20417 12851 20451
rect 13645 20417 13679 20451
rect 13912 20417 13946 20451
rect 17969 20417 18003 20451
rect 19901 20417 19935 20451
rect 21833 20417 21867 20451
rect 23121 20417 23155 20451
rect 23388 20417 23422 20451
rect 24961 20417 24995 20451
rect 26433 20417 26467 20451
rect 27353 20417 27387 20451
rect 27445 20417 27479 20451
rect 28641 20417 28675 20451
rect 29009 20417 29043 20451
rect 30297 20417 30331 20451
rect 31401 20417 31435 20451
rect 32781 20417 32815 20451
rect 33517 20417 33551 20451
rect 16681 20349 16715 20383
rect 16957 20349 16991 20383
rect 21005 20349 21039 20383
rect 21189 20349 21223 20383
rect 25237 20349 25271 20383
rect 26985 20349 27019 20383
rect 27169 20349 27203 20383
rect 27261 20349 27295 20383
rect 28733 20349 28767 20383
rect 29101 20349 29135 20383
rect 30389 20349 30423 20383
rect 30481 20349 30515 20383
rect 32873 20349 32907 20383
rect 19349 20281 19383 20315
rect 29929 20281 29963 20315
rect 16037 20213 16071 20247
rect 20545 20213 20579 20247
rect 22201 20213 22235 20247
rect 24501 20213 24535 20247
rect 31493 20213 31527 20247
rect 13369 20009 13403 20043
rect 19809 20009 19843 20043
rect 21925 20009 21959 20043
rect 23397 20009 23431 20043
rect 26341 20009 26375 20043
rect 27721 20009 27755 20043
rect 30573 20009 30607 20043
rect 32413 20009 32447 20043
rect 20821 19941 20855 19975
rect 23765 19941 23799 19975
rect 24869 19941 24903 19975
rect 27629 19941 27663 19975
rect 35357 19941 35391 19975
rect 17877 19873 17911 19907
rect 20177 19873 20211 19907
rect 22293 19873 22327 19907
rect 28457 19873 28491 19907
rect 31125 19873 31159 19907
rect 32965 19873 32999 19907
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 15025 19805 15059 19839
rect 15669 19805 15703 19839
rect 17509 19805 17543 19839
rect 17693 19805 17727 19839
rect 17785 19805 17819 19839
rect 18061 19805 18095 19839
rect 19993 19805 20027 19839
rect 20085 19805 20119 19839
rect 20269 19805 20303 19839
rect 21097 19805 21131 19839
rect 21202 19799 21236 19833
rect 21302 19805 21336 19839
rect 21465 19805 21499 19839
rect 22109 19805 22143 19839
rect 22201 19805 22235 19839
rect 22385 19805 22419 19839
rect 23581 19805 23615 19839
rect 23857 19805 23891 19839
rect 24593 19805 24627 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 25053 19805 25087 19839
rect 25973 19805 26007 19839
rect 26341 19805 26375 19839
rect 29929 19805 29963 19839
rect 30941 19805 30975 19839
rect 31769 19805 31803 19839
rect 32781 19805 32815 19839
rect 33609 19805 33643 19839
rect 35173 19805 35207 19839
rect 14473 19737 14507 19771
rect 15209 19737 15243 19771
rect 15936 19737 15970 19771
rect 27261 19737 27295 19771
rect 28273 19737 28307 19771
rect 32873 19737 32907 19771
rect 17049 19669 17083 19703
rect 18245 19669 18279 19703
rect 26525 19669 26559 19703
rect 30021 19669 30055 19703
rect 31033 19669 31067 19703
rect 31861 19669 31895 19703
rect 33701 19669 33735 19703
rect 19441 19465 19475 19499
rect 21189 19465 21223 19499
rect 24777 19465 24811 19499
rect 26985 19465 27019 19499
rect 27445 19465 27479 19499
rect 28089 19465 28123 19499
rect 32505 19465 32539 19499
rect 32965 19465 32999 19499
rect 33793 19465 33827 19499
rect 13461 19397 13495 19431
rect 14749 19397 14783 19431
rect 20913 19397 20947 19431
rect 21925 19397 21959 19431
rect 30205 19397 30239 19431
rect 32873 19397 32907 19431
rect 12265 19329 12299 19363
rect 15485 19329 15519 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17233 19329 17267 19363
rect 18337 19329 18371 19363
rect 18521 19329 18555 19363
rect 19717 19329 19751 19363
rect 19809 19329 19843 19363
rect 19901 19329 19935 19363
rect 20085 19329 20119 19363
rect 20545 19329 20579 19363
rect 20638 19329 20672 19363
rect 20821 19329 20855 19363
rect 21051 19329 21085 19363
rect 22836 19329 22870 19363
rect 24685 19329 24719 19363
rect 25421 19329 25455 19363
rect 27537 19329 27571 19363
rect 28343 19329 28377 19363
rect 29377 19329 29411 19363
rect 29561 19329 29595 19363
rect 30849 19329 30883 19363
rect 33701 19329 33735 19363
rect 28549 19295 28583 19329
rect 16957 19261 16991 19295
rect 18153 19261 18187 19295
rect 18613 19261 18647 19295
rect 22109 19261 22143 19295
rect 22569 19261 22603 19295
rect 25697 19261 25731 19295
rect 27169 19261 27203 19295
rect 27261 19261 27295 19295
rect 27629 19261 27663 19295
rect 28265 19261 28299 19295
rect 28457 19261 28491 19295
rect 29653 19261 29687 19295
rect 33149 19261 33183 19295
rect 14933 19193 14967 19227
rect 30389 19193 30423 19227
rect 12081 19125 12115 19159
rect 13553 19125 13587 19159
rect 15577 19125 15611 19159
rect 17417 19125 17451 19159
rect 23949 19125 23983 19159
rect 29193 19125 29227 19159
rect 30941 19125 30975 19159
rect 13461 18921 13495 18955
rect 16405 18921 16439 18955
rect 20085 18921 20119 18955
rect 21189 18921 21223 18955
rect 23305 18921 23339 18955
rect 27445 18921 27479 18955
rect 30021 18921 30055 18955
rect 31125 18921 31159 18955
rect 32137 18921 32171 18955
rect 33885 18921 33919 18955
rect 22293 18853 22327 18887
rect 23581 18853 23615 18887
rect 23673 18853 23707 18887
rect 16865 18785 16899 18819
rect 17785 18785 17819 18819
rect 17877 18785 17911 18819
rect 25329 18785 25363 18819
rect 25605 18785 25639 18819
rect 27629 18785 27663 18819
rect 27813 18785 27847 18819
rect 32321 18785 32355 18819
rect 11437 18717 11471 18751
rect 14105 18717 14139 18751
rect 16589 18717 16623 18751
rect 16773 18717 16807 18751
rect 17509 18717 17543 18751
rect 17693 18717 17727 18751
rect 18061 18717 18095 18751
rect 19441 18717 19475 18751
rect 19534 18717 19568 18751
rect 19717 18717 19751 18751
rect 19947 18717 19981 18751
rect 20545 18717 20579 18751
rect 20638 18717 20672 18751
rect 20821 18717 20855 18751
rect 21010 18717 21044 18751
rect 21649 18717 21683 18751
rect 21742 18717 21776 18751
rect 21925 18717 21959 18751
rect 22155 18717 22189 18751
rect 23489 18717 23523 18751
rect 23765 18717 23799 18751
rect 24777 18717 24811 18751
rect 26985 18717 27019 18751
rect 27721 18717 27755 18751
rect 27905 18717 27939 18751
rect 28457 18717 28491 18751
rect 28733 18717 28767 18751
rect 28825 18717 28859 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 30481 18717 30515 18751
rect 30573 18717 30607 18751
rect 31033 18717 31067 18751
rect 31861 18717 31895 18751
rect 32781 18717 32815 18751
rect 33057 18717 33091 18751
rect 33149 18717 33183 18751
rect 33793 18717 33827 18751
rect 11682 18649 11716 18683
rect 13369 18649 13403 18683
rect 14350 18649 14384 18683
rect 19809 18649 19843 18683
rect 20913 18649 20947 18683
rect 22014 18649 22048 18683
rect 24593 18649 24627 18683
rect 25053 18649 25087 18683
rect 28641 18649 28675 18683
rect 32965 18649 32999 18683
rect 12817 18581 12851 18615
rect 15485 18581 15519 18615
rect 18245 18581 18279 18615
rect 24961 18581 24995 18615
rect 26525 18581 26559 18615
rect 26801 18581 26835 18615
rect 29009 18581 29043 18615
rect 33333 18581 33367 18615
rect 15117 18377 15151 18411
rect 21281 18377 21315 18411
rect 22109 18377 22143 18411
rect 27353 18377 27387 18411
rect 29193 18377 29227 18411
rect 30389 18377 30423 18411
rect 21005 18309 21039 18343
rect 25145 18309 25179 18343
rect 26433 18309 26467 18343
rect 31033 18309 31067 18343
rect 33977 18309 34011 18343
rect 11785 18241 11819 18275
rect 13737 18241 13771 18275
rect 14004 18241 14038 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 17969 18241 18003 18275
rect 18236 18241 18270 18275
rect 20177 18241 20211 18275
rect 20637 18241 20671 18275
rect 20730 18241 20764 18275
rect 20913 18241 20947 18275
rect 21143 18241 21177 18275
rect 22385 18241 22419 18275
rect 22474 18247 22508 18281
rect 22569 18241 22603 18275
rect 22753 18241 22787 18275
rect 23581 18241 23615 18275
rect 24317 18241 24351 18275
rect 24409 18241 24443 18275
rect 24501 18241 24535 18275
rect 24685 18241 24719 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 26249 18241 26283 18275
rect 27169 18241 27203 18275
rect 27261 18241 27295 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 28549 18241 28583 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 29929 18241 29963 18275
rect 30665 18241 30699 18275
rect 30941 18241 30975 18275
rect 32965 18241 32999 18275
rect 33057 18241 33091 18275
rect 33333 18241 33367 18275
rect 33793 18241 33827 18275
rect 34069 18241 34103 18275
rect 34166 18247 34200 18281
rect 11529 18173 11563 18207
rect 16129 18173 16163 18207
rect 16865 18173 16899 18207
rect 17141 18173 17175 18207
rect 19625 18173 19659 18207
rect 27537 18173 27571 18207
rect 28273 18173 28307 18207
rect 28365 18173 28399 18207
rect 30573 18173 30607 18207
rect 25145 18105 25179 18139
rect 29469 18105 29503 18139
rect 29653 18105 29687 18139
rect 33793 18105 33827 18139
rect 12909 18037 12943 18071
rect 15669 18037 15703 18071
rect 19349 18037 19383 18071
rect 19993 18037 20027 18071
rect 23029 18037 23063 18071
rect 23397 18037 23431 18071
rect 24041 18037 24075 18071
rect 27445 18037 27479 18071
rect 28733 18037 28767 18071
rect 32781 18037 32815 18071
rect 33241 18037 33275 18071
rect 10793 17833 10827 17867
rect 14565 17833 14599 17867
rect 17049 17833 17083 17867
rect 18245 17833 18279 17867
rect 19257 17833 19291 17867
rect 21189 17833 21223 17867
rect 22201 17833 22235 17867
rect 28181 17833 28215 17867
rect 28825 17833 28859 17867
rect 29929 17833 29963 17867
rect 19625 17765 19659 17799
rect 28917 17765 28951 17799
rect 30665 17765 30699 17799
rect 31493 17765 31527 17799
rect 33241 17765 33275 17799
rect 11437 17697 11471 17731
rect 13553 17697 13587 17731
rect 15025 17697 15059 17731
rect 17877 17697 17911 17731
rect 26801 17697 26835 17731
rect 29009 17697 29043 17731
rect 31769 17697 31803 17731
rect 32229 17697 32263 17731
rect 32689 17697 32723 17731
rect 11704 17629 11738 17663
rect 13369 17629 13403 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 15669 17629 15703 17663
rect 15936 17629 15970 17663
rect 17509 17629 17543 17663
rect 17693 17629 17727 17663
rect 17785 17629 17819 17663
rect 18061 17629 18095 17663
rect 19441 17629 19475 17663
rect 19717 17629 19751 17663
rect 20545 17629 20579 17663
rect 20638 17629 20672 17663
rect 20821 17629 20855 17663
rect 21010 17629 21044 17663
rect 22937 17629 22971 17663
rect 23029 17629 23063 17663
rect 23121 17629 23155 17663
rect 23305 17629 23339 17663
rect 24869 17629 24903 17663
rect 27057 17629 27091 17663
rect 28733 17629 28767 17663
rect 29561 17629 29595 17663
rect 29929 17629 29963 17663
rect 30113 17629 30147 17663
rect 30665 17629 30699 17663
rect 30849 17629 30883 17663
rect 31401 17629 31435 17663
rect 32413 17629 32447 17663
rect 32505 17629 32539 17663
rect 32781 17629 32815 17663
rect 33614 17629 33648 17663
rect 10609 17561 10643 17595
rect 10825 17561 10859 17595
rect 20913 17561 20947 17595
rect 21833 17561 21867 17595
rect 22017 17561 22051 17595
rect 25114 17561 25148 17595
rect 31493 17561 31527 17595
rect 33241 17561 33275 17595
rect 33425 17561 33459 17595
rect 33517 17561 33551 17595
rect 10977 17493 11011 17527
rect 12817 17493 12851 17527
rect 22661 17493 22695 17527
rect 26249 17493 26283 17527
rect 29745 17493 29779 17527
rect 31585 17493 31619 17527
rect 11897 17289 11931 17323
rect 12567 17289 12601 17323
rect 13645 17289 13679 17323
rect 15301 17289 15335 17323
rect 16129 17289 16163 17323
rect 24593 17289 24627 17323
rect 25973 17289 26007 17323
rect 28457 17289 28491 17323
rect 29193 17289 29227 17323
rect 31585 17289 31619 17323
rect 32597 17289 32631 17323
rect 11529 17221 11563 17255
rect 11745 17221 11779 17255
rect 12403 17221 12437 17255
rect 16773 17221 16807 17255
rect 17938 17221 17972 17255
rect 22998 17221 23032 17255
rect 10977 17153 11011 17187
rect 13829 17153 13863 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 15117 17153 15151 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16957 17153 16991 17187
rect 17141 17153 17175 17187
rect 17233 17153 17267 17187
rect 19533 17153 19567 17187
rect 22047 17153 22081 17187
rect 24869 17153 24903 17187
rect 24961 17153 24995 17187
rect 25053 17153 25087 17187
rect 25237 17153 25271 17187
rect 25881 17153 25915 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 28089 17153 28123 17187
rect 29377 17153 29411 17187
rect 30113 17153 30147 17187
rect 30481 17153 30515 17187
rect 31217 17153 31251 17187
rect 31309 17153 31343 17187
rect 31401 17153 31435 17187
rect 32229 17153 32263 17187
rect 32321 17153 32355 17187
rect 32413 17153 32447 17187
rect 14105 17085 14139 17119
rect 14841 17085 14875 17119
rect 14933 17085 14967 17119
rect 17693 17085 17727 17119
rect 22293 17085 22327 17119
rect 22753 17085 22787 17119
rect 28181 17085 28215 17119
rect 29653 17085 29687 17119
rect 10793 17017 10827 17051
rect 12725 17017 12759 17051
rect 19073 17017 19107 17051
rect 29561 17017 29595 17051
rect 30665 17017 30699 17051
rect 11713 16949 11747 16983
rect 12541 16949 12575 16983
rect 14013 16949 14047 16983
rect 20821 16949 20855 16983
rect 21833 16949 21867 16983
rect 22201 16949 22235 16983
rect 24133 16949 24167 16983
rect 27077 16949 27111 16983
rect 28273 16949 28307 16983
rect 30389 16949 30423 16983
rect 12173 16745 12207 16779
rect 15025 16745 15059 16779
rect 18429 16745 18463 16779
rect 19993 16745 20027 16779
rect 20913 16745 20947 16779
rect 21465 16745 21499 16779
rect 28549 16745 28583 16779
rect 30297 16745 30331 16779
rect 33977 16745 34011 16779
rect 17233 16677 17267 16711
rect 27261 16677 27295 16711
rect 11529 16609 11563 16643
rect 14565 16609 14599 16643
rect 16405 16609 16439 16643
rect 17969 16609 18003 16643
rect 19625 16609 19659 16643
rect 20729 16609 20763 16643
rect 21925 16609 21959 16643
rect 25881 16609 25915 16643
rect 31401 16609 31435 16643
rect 32873 16609 32907 16643
rect 10793 16541 10827 16575
rect 11345 16541 11379 16575
rect 12725 16541 12759 16575
rect 13001 16541 13035 16575
rect 14289 16541 14323 16575
rect 14473 16541 14507 16575
rect 14657 16541 14691 16575
rect 14841 16541 14875 16575
rect 15669 16541 15703 16575
rect 16865 16541 16899 16575
rect 17049 16541 17083 16575
rect 17693 16541 17727 16575
rect 17877 16541 17911 16575
rect 18061 16541 18095 16575
rect 18245 16541 18279 16575
rect 19257 16541 19291 16575
rect 19441 16541 19475 16575
rect 19533 16541 19567 16575
rect 19809 16541 19843 16575
rect 20637 16541 20671 16575
rect 21649 16541 21683 16575
rect 21833 16541 21867 16575
rect 23075 16541 23109 16575
rect 23213 16541 23247 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 25033 16541 25067 16575
rect 25145 16541 25179 16575
rect 25237 16541 25271 16575
rect 25421 16541 25455 16575
rect 27721 16541 27755 16575
rect 27905 16541 27939 16575
rect 28457 16541 28491 16575
rect 31125 16541 31159 16575
rect 32413 16541 32447 16575
rect 32781 16541 32815 16575
rect 32965 16541 32999 16575
rect 33609 16541 33643 16575
rect 33701 16541 33735 16575
rect 33793 16541 33827 16575
rect 12081 16473 12115 16507
rect 16221 16473 16255 16507
rect 21005 16473 21039 16507
rect 22845 16473 22879 16507
rect 26126 16473 26160 16507
rect 30205 16473 30239 16507
rect 10609 16405 10643 16439
rect 15485 16405 15519 16439
rect 24777 16405 24811 16439
rect 27905 16405 27939 16439
rect 22201 16201 22235 16235
rect 26341 16201 26375 16235
rect 30297 16201 30331 16235
rect 32689 16201 32723 16235
rect 33333 16201 33367 16235
rect 13369 16133 13403 16167
rect 13569 16133 13603 16167
rect 22017 16133 22051 16167
rect 26157 16133 26191 16167
rect 10425 16065 10459 16099
rect 12173 16065 12207 16099
rect 12725 16065 12759 16099
rect 12909 16065 12943 16099
rect 14473 16065 14507 16099
rect 14657 16065 14691 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 15853 16065 15887 16099
rect 16681 16065 16715 16099
rect 16957 16065 16991 16099
rect 18613 16065 18647 16099
rect 19809 16065 19843 16099
rect 20076 16065 20110 16099
rect 21833 16065 21867 16099
rect 24133 16065 24167 16099
rect 24400 16065 24434 16099
rect 25973 16065 26007 16099
rect 27077 16065 27111 16099
rect 27997 16065 28031 16099
rect 28089 16065 28123 16099
rect 28181 16065 28215 16099
rect 28365 16065 28399 16099
rect 28825 16065 28859 16099
rect 29745 16065 29779 16099
rect 30113 16065 30147 16099
rect 30757 16065 30791 16099
rect 32137 16065 32171 16099
rect 33241 16065 33275 16099
rect 14749 15997 14783 16031
rect 14841 15997 14875 16031
rect 16129 15997 16163 16031
rect 18337 15997 18371 16031
rect 22845 15997 22879 16031
rect 23121 15997 23155 16031
rect 31033 15997 31067 16031
rect 32413 15997 32447 16031
rect 13737 15929 13771 15963
rect 27169 15929 27203 15963
rect 10241 15861 10275 15895
rect 11989 15861 12023 15895
rect 13553 15861 13587 15895
rect 15669 15861 15703 15895
rect 16037 15861 16071 15895
rect 21189 15861 21223 15895
rect 25513 15861 25547 15895
rect 27721 15861 27755 15895
rect 28917 15861 28951 15895
rect 30113 15861 30147 15895
rect 32505 15861 32539 15895
rect 13553 15657 13587 15691
rect 18521 15657 18555 15691
rect 24409 15657 24443 15691
rect 30941 15657 30975 15691
rect 10885 15589 10919 15623
rect 21189 15589 21223 15623
rect 26893 15589 26927 15623
rect 11713 15521 11747 15555
rect 15025 15521 15059 15555
rect 16313 15521 16347 15555
rect 17049 15521 17083 15555
rect 17325 15521 17359 15555
rect 19257 15521 19291 15555
rect 21649 15521 21683 15555
rect 21741 15521 21775 15555
rect 25513 15521 25547 15555
rect 29561 15521 29595 15555
rect 31677 15521 31711 15555
rect 9505 15453 9539 15487
rect 12173 15453 12207 15487
rect 12429 15453 12463 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 14933 15453 14967 15487
rect 15209 15453 15243 15487
rect 16037 15453 16071 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 16589 15453 16623 15487
rect 18245 15453 18279 15487
rect 18705 15453 18739 15487
rect 19533 15453 19567 15487
rect 20545 15453 20579 15487
rect 22661 15453 22695 15487
rect 22937 15453 22971 15487
rect 24685 15453 24719 15487
rect 24774 15453 24808 15487
rect 24869 15453 24903 15487
rect 25053 15453 25087 15487
rect 25769 15453 25803 15487
rect 28089 15453 28123 15487
rect 28181 15453 28215 15487
rect 28273 15453 28307 15487
rect 28457 15453 28491 15487
rect 29817 15453 29851 15487
rect 31401 15453 31435 15487
rect 9772 15385 9806 15419
rect 11345 15385 11379 15419
rect 11529 15385 11563 15419
rect 20637 15385 20671 15419
rect 15393 15317 15427 15351
rect 16773 15317 16807 15351
rect 21557 15317 21591 15351
rect 27813 15317 27847 15351
rect 8861 15113 8895 15147
rect 21833 15113 21867 15147
rect 26433 15113 26467 15147
rect 30665 15113 30699 15147
rect 31309 15113 31343 15147
rect 9772 15045 9806 15079
rect 27353 15045 27387 15079
rect 31217 15045 31251 15079
rect 9045 14977 9079 15011
rect 9505 14977 9539 15011
rect 12081 14977 12115 15011
rect 12348 14977 12382 15011
rect 14648 14977 14682 15011
rect 16865 14977 16899 15011
rect 17141 14977 17175 15011
rect 18153 14977 18187 15011
rect 18889 14977 18923 15011
rect 19073 14977 19107 15011
rect 19257 14977 19291 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 21189 14977 21223 15011
rect 22017 14977 22051 15011
rect 22477 14977 22511 15011
rect 24225 14977 24259 15011
rect 24314 14983 24348 15017
rect 24409 14980 24443 15014
rect 24593 14977 24627 15011
rect 25053 14977 25087 15011
rect 25309 14977 25343 15011
rect 26985 14977 27019 15011
rect 27169 14977 27203 15011
rect 28089 14977 28123 15011
rect 28181 14977 28215 15011
rect 28273 14977 28307 15011
rect 28457 14977 28491 15011
rect 29285 14977 29319 15011
rect 29541 14977 29575 15011
rect 14381 14909 14415 14943
rect 19159 14909 19193 14943
rect 20545 14909 20579 14943
rect 23949 14909 23983 14943
rect 15761 14841 15795 14875
rect 20085 14841 20119 14875
rect 22845 14841 22879 14875
rect 10885 14773 10919 14807
rect 13461 14773 13495 14807
rect 18337 14773 18371 14807
rect 21005 14773 21039 14807
rect 22937 14773 22971 14807
rect 27813 14773 27847 14807
rect 13093 14569 13127 14603
rect 15669 14569 15703 14603
rect 17509 14569 17543 14603
rect 21373 14569 21407 14603
rect 25697 14569 25731 14603
rect 26709 14569 26743 14603
rect 28825 14569 28859 14603
rect 30941 14569 30975 14603
rect 12173 14501 12207 14535
rect 25881 14501 25915 14535
rect 9505 14433 9539 14467
rect 18337 14433 18371 14467
rect 19993 14433 20027 14467
rect 29561 14433 29595 14467
rect 9772 14365 9806 14399
rect 11713 14365 11747 14399
rect 12357 14365 12391 14399
rect 14289 14365 14323 14399
rect 16129 14365 16163 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 18245 14365 18279 14399
rect 18521 14365 18555 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 22661 14365 22695 14399
rect 22754 14365 22788 14399
rect 23126 14365 23160 14399
rect 24409 14365 24443 14399
rect 24502 14365 24536 14399
rect 24685 14365 24719 14399
rect 24874 14365 24908 14399
rect 27445 14365 27479 14399
rect 27629 14365 27663 14399
rect 28273 14365 28307 14399
rect 28733 14365 28767 14399
rect 28917 14365 28951 14399
rect 29817 14365 29851 14399
rect 11345 14297 11379 14331
rect 11529 14297 11563 14331
rect 12909 14297 12943 14331
rect 13125 14297 13159 14331
rect 14556 14297 14590 14331
rect 16396 14297 16430 14331
rect 19349 14297 19383 14331
rect 20260 14297 20294 14331
rect 22937 14297 22971 14331
rect 23029 14297 23063 14331
rect 24777 14297 24811 14331
rect 25513 14297 25547 14331
rect 26525 14297 26559 14331
rect 10885 14229 10919 14263
rect 13277 14229 13311 14263
rect 18705 14229 18739 14263
rect 19441 14229 19475 14263
rect 22201 14229 22235 14263
rect 23305 14229 23339 14263
rect 25053 14229 25087 14263
rect 25713 14229 25747 14263
rect 26725 14229 26759 14263
rect 26893 14229 26927 14263
rect 28089 14229 28123 14263
rect 8861 14025 8895 14059
rect 10885 14025 10919 14059
rect 12725 14025 12759 14059
rect 13185 14025 13219 14059
rect 14933 14025 14967 14059
rect 16681 14025 16715 14059
rect 22661 14025 22695 14059
rect 24593 14025 24627 14059
rect 28549 14025 28583 14059
rect 29745 14025 29779 14059
rect 11713 13957 11747 13991
rect 12541 13957 12575 13991
rect 16129 13957 16163 13991
rect 26065 13957 26099 13991
rect 26265 13957 26299 13991
rect 9045 13889 9079 13923
rect 9772 13889 9806 13923
rect 11529 13889 11563 13923
rect 12357 13889 12391 13923
rect 13369 13889 13403 13923
rect 14473 13889 14507 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 15945 13889 15979 13923
rect 16865 13889 16899 13923
rect 17141 13889 17175 13923
rect 18061 13889 18095 13923
rect 18245 13889 18279 13923
rect 18429 13889 18463 13923
rect 18613 13889 18647 13923
rect 19257 13889 19291 13923
rect 19441 13895 19475 13929
rect 19533 13889 19567 13923
rect 19809 13889 19843 13923
rect 20637 13889 20671 13923
rect 20821 13889 20855 13923
rect 21833 13889 21867 13923
rect 22017 13889 22051 13923
rect 22845 13889 22879 13923
rect 24777 13889 24811 13923
rect 24869 13889 24903 13923
rect 25145 13889 25179 13923
rect 27169 13889 27203 13923
rect 27436 13889 27470 13923
rect 29193 13889 29227 13923
rect 29653 13889 29687 13923
rect 29837 13889 29871 13923
rect 9505 13821 9539 13855
rect 15393 13821 15427 13855
rect 17049 13821 17083 13855
rect 18337 13821 18371 13855
rect 19625 13821 19659 13855
rect 20913 13821 20947 13855
rect 22201 13821 22235 13855
rect 23305 13821 23339 13855
rect 23581 13821 23615 13855
rect 20453 13753 20487 13787
rect 25053 13753 25087 13787
rect 11897 13685 11931 13719
rect 14289 13685 14323 13719
rect 18797 13685 18831 13719
rect 19993 13685 20027 13719
rect 26249 13685 26283 13719
rect 26433 13685 26467 13719
rect 29009 13685 29043 13719
rect 10885 13481 10919 13515
rect 11713 13481 11747 13515
rect 21097 13481 21131 13515
rect 25697 13481 25731 13515
rect 28181 13481 28215 13515
rect 13369 13413 13403 13447
rect 17233 13413 17267 13447
rect 25053 13413 25087 13447
rect 29009 13413 29043 13447
rect 19717 13345 19751 13379
rect 23213 13345 23247 13379
rect 23305 13345 23339 13379
rect 9505 13277 9539 13311
rect 9772 13277 9806 13311
rect 11529 13277 11563 13311
rect 12265 13277 12299 13311
rect 13185 13277 13219 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 14933 13277 14967 13311
rect 15577 13277 15611 13311
rect 16221 13277 16255 13311
rect 17049 13277 17083 13311
rect 18429 13277 18463 13311
rect 18613 13277 18647 13311
rect 18705 13277 18739 13311
rect 22201 13277 22235 13311
rect 22477 13277 22511 13311
rect 23121 13277 23155 13311
rect 23397 13277 23431 13311
rect 23581 13277 23615 13311
rect 24409 13277 24443 13311
rect 24502 13277 24536 13311
rect 24685 13277 24719 13311
rect 24777 13277 24811 13311
rect 24874 13277 24908 13311
rect 25513 13277 25547 13311
rect 26709 13277 26743 13311
rect 26857 13277 26891 13311
rect 27215 13277 27249 13311
rect 28641 13277 28675 13311
rect 28825 13277 28859 13311
rect 11345 13209 11379 13243
rect 12449 13209 12483 13243
rect 14197 13209 14231 13243
rect 19984 13209 20018 13243
rect 22017 13209 22051 13243
rect 26985 13209 27019 13243
rect 27077 13209 27111 13243
rect 27813 13209 27847 13243
rect 27997 13209 28031 13243
rect 12633 13141 12667 13175
rect 14749 13141 14783 13175
rect 15393 13141 15427 13175
rect 16037 13141 16071 13175
rect 18245 13141 18279 13175
rect 22385 13141 22419 13175
rect 22937 13141 22971 13175
rect 27353 13141 27387 13175
rect 10241 12937 10275 12971
rect 13001 12937 13035 12971
rect 14841 12937 14875 12971
rect 20085 12937 20119 12971
rect 25237 12937 25271 12971
rect 30021 12937 30055 12971
rect 11888 12869 11922 12903
rect 13728 12869 13762 12903
rect 18398 12869 18432 12903
rect 24961 12869 24995 12903
rect 25697 12869 25731 12903
rect 25897 12869 25931 12903
rect 27261 12869 27295 12903
rect 27353 12869 27387 12903
rect 28908 12869 28942 12903
rect 9781 12801 9815 12835
rect 10425 12801 10459 12835
rect 13461 12801 13495 12835
rect 15485 12801 15519 12835
rect 16129 12801 16163 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 17693 12801 17727 12835
rect 20269 12801 20303 12835
rect 20453 12801 20487 12835
rect 21097 12801 21131 12835
rect 21281 12801 21315 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 23020 12801 23054 12835
rect 24593 12801 24627 12835
rect 24686 12801 24720 12835
rect 24869 12801 24903 12835
rect 25058 12801 25092 12835
rect 26985 12801 27019 12835
rect 27078 12801 27112 12835
rect 27450 12801 27484 12835
rect 28641 12801 28675 12835
rect 11621 12733 11655 12767
rect 16681 12733 16715 12767
rect 18153 12733 18187 12767
rect 20545 12733 20579 12767
rect 22753 12733 22787 12767
rect 9597 12665 9631 12699
rect 15945 12665 15979 12699
rect 19533 12665 19567 12699
rect 24133 12665 24167 12699
rect 15301 12597 15335 12631
rect 17509 12597 17543 12631
rect 21097 12597 21131 12631
rect 22201 12597 22235 12631
rect 25881 12597 25915 12631
rect 26065 12597 26099 12631
rect 27629 12597 27663 12631
rect 11805 12393 11839 12427
rect 12449 12393 12483 12427
rect 14473 12393 14507 12427
rect 17601 12393 17635 12427
rect 25329 12393 25363 12427
rect 20637 12325 20671 12359
rect 22569 12325 22603 12359
rect 23489 12325 23523 12359
rect 14105 12257 14139 12291
rect 16221 12257 16255 12291
rect 27629 12257 27663 12291
rect 9137 12189 9171 12223
rect 10241 12189 10275 12223
rect 10885 12189 10919 12223
rect 11989 12189 12023 12223
rect 12633 12189 12667 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 14933 12189 14967 12223
rect 15301 12189 15335 12223
rect 16488 12189 16522 12223
rect 18245 12189 18279 12223
rect 19257 12189 19291 12223
rect 21189 12189 21223 12223
rect 23213 12189 23247 12223
rect 23305 12189 23339 12223
rect 23581 12189 23615 12223
rect 24685 12189 24719 12223
rect 26157 12189 26191 12223
rect 26250 12189 26284 12223
rect 26433 12189 26467 12223
rect 26663 12189 26697 12223
rect 29745 12189 29779 12223
rect 15117 12121 15151 12155
rect 15209 12121 15243 12155
rect 19524 12121 19558 12155
rect 21434 12121 21468 12155
rect 25145 12121 25179 12155
rect 26525 12121 26559 12155
rect 27896 12121 27930 12155
rect 8953 12053 8987 12087
rect 10057 12053 10091 12087
rect 10701 12053 10735 12087
rect 13369 12053 13403 12087
rect 15485 12053 15519 12087
rect 18061 12053 18095 12087
rect 23029 12053 23063 12087
rect 24501 12053 24535 12087
rect 25345 12053 25379 12087
rect 25513 12053 25547 12087
rect 26801 12053 26835 12087
rect 29009 12053 29043 12087
rect 29561 12053 29595 12087
rect 11897 11849 11931 11883
rect 14105 11849 14139 11883
rect 15945 11849 15979 11883
rect 20269 11849 20303 11883
rect 21281 11849 21315 11883
rect 23489 11849 23523 11883
rect 25989 11849 26023 11883
rect 27997 11849 28031 11883
rect 29929 11849 29963 11883
rect 9658 11781 9692 11815
rect 17224 11781 17258 11815
rect 20913 11781 20947 11815
rect 24159 11781 24193 11815
rect 24333 11781 24367 11815
rect 24961 11781 24995 11815
rect 25177 11781 25211 11815
rect 25789 11781 25823 11815
rect 27629 11781 27663 11815
rect 28816 11781 28850 11815
rect 21143 11747 21177 11781
rect 7748 11713 7782 11747
rect 11713 11713 11747 11747
rect 12725 11713 12759 11747
rect 12992 11713 13026 11747
rect 14565 11713 14599 11747
rect 14832 11713 14866 11747
rect 16957 11713 16991 11747
rect 18981 11713 19015 11747
rect 19625 11713 19659 11747
rect 20453 11713 20487 11747
rect 22385 11713 22419 11747
rect 23397 11713 23431 11747
rect 23581 11713 23615 11747
rect 27169 11713 27203 11747
rect 27813 11713 27847 11747
rect 28549 11713 28583 11747
rect 7481 11645 7515 11679
rect 9413 11645 9447 11679
rect 11529 11645 11563 11679
rect 22109 11645 22143 11679
rect 25329 11577 25363 11611
rect 26985 11577 27019 11611
rect 8861 11509 8895 11543
rect 10793 11509 10827 11543
rect 18337 11509 18371 11543
rect 18797 11509 18831 11543
rect 19441 11509 19475 11543
rect 21097 11509 21131 11543
rect 24317 11509 24351 11543
rect 24501 11509 24535 11543
rect 25145 11509 25179 11543
rect 25973 11509 26007 11543
rect 26157 11509 26191 11543
rect 8953 11305 8987 11339
rect 14749 11305 14783 11339
rect 16773 11305 16807 11339
rect 24685 11305 24719 11339
rect 28457 11305 28491 11339
rect 30205 11305 30239 11339
rect 31493 11305 31527 11339
rect 7941 11237 7975 11271
rect 13001 11237 13035 11271
rect 15761 11237 15795 11271
rect 20637 11237 20671 11271
rect 27169 11237 27203 11271
rect 19257 11169 19291 11203
rect 21741 11169 21775 11203
rect 23581 11169 23615 11203
rect 6561 11101 6595 11135
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 11621 11101 11655 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 15209 11101 15243 11135
rect 15577 11101 15611 11135
rect 16221 11101 16255 11135
rect 16497 11101 16531 11135
rect 16613 11101 16647 11135
rect 17253 11101 17287 11135
rect 17509 11101 17543 11135
rect 17601 11101 17635 11135
rect 18429 11101 18463 11135
rect 21281 11101 21315 11135
rect 21373 11101 21407 11135
rect 21557 11101 21591 11135
rect 22753 11101 22787 11135
rect 23489 11101 23523 11135
rect 23673 11101 23707 11135
rect 25421 11101 25455 11135
rect 25514 11101 25548 11135
rect 25697 11101 25731 11135
rect 25886 11101 25920 11135
rect 26525 11101 26559 11135
rect 26618 11101 26652 11135
rect 26990 11101 27024 11135
rect 27629 11101 27663 11135
rect 27813 11101 27847 11135
rect 27997 11101 28031 11135
rect 28641 11101 28675 11135
rect 29745 11101 29779 11135
rect 30389 11101 30423 11135
rect 31033 11101 31067 11135
rect 31677 11101 31711 11135
rect 6806 11033 6840 11067
rect 10048 11033 10082 11067
rect 11866 11033 11900 11067
rect 15393 11033 15427 11067
rect 15485 11033 15519 11067
rect 16405 11033 16439 11067
rect 17417 11033 17451 11067
rect 19502 11033 19536 11067
rect 24593 11033 24627 11067
rect 25789 11033 25823 11067
rect 26801 11033 26835 11067
rect 26893 11033 26927 11067
rect 11161 10965 11195 10999
rect 17785 10965 17819 10999
rect 18245 10965 18279 10999
rect 22937 10965 22971 10999
rect 26065 10965 26099 10999
rect 29561 10965 29595 10999
rect 30849 10965 30883 10999
rect 6469 10761 6503 10795
rect 7481 10761 7515 10795
rect 10977 10761 11011 10795
rect 11897 10761 11931 10795
rect 14105 10761 14139 10795
rect 17141 10761 17175 10795
rect 19901 10761 19935 10795
rect 29101 10761 29135 10795
rect 15301 10693 15335 10727
rect 15393 10693 15427 10727
rect 23673 10693 23707 10727
rect 30297 10693 30331 10727
rect 6653 10625 6687 10659
rect 7297 10625 7331 10659
rect 8125 10625 8159 10659
rect 8953 10625 8987 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 13921 10625 13955 10659
rect 15117 10625 15151 10659
rect 15485 10625 15519 10659
rect 16957 10625 16991 10659
rect 17785 10625 17819 10659
rect 18797 10625 18831 10659
rect 19441 10625 19475 10659
rect 19717 10625 19751 10659
rect 20637 10625 20671 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 21833 10625 21867 10659
rect 22753 10625 22787 10659
rect 23397 10625 23431 10659
rect 23490 10625 23524 10659
rect 23765 10625 23799 10659
rect 23903 10625 23937 10659
rect 24869 10625 24903 10659
rect 25881 10625 25915 10659
rect 27077 10625 27111 10659
rect 27721 10625 27755 10659
rect 27988 10625 28022 10659
rect 30113 10625 30147 10659
rect 30941 10625 30975 10659
rect 31585 10625 31619 10659
rect 7113 10557 7147 10591
rect 10609 10557 10643 10591
rect 12449 10557 12483 10591
rect 12725 10557 12759 10591
rect 13737 10557 13771 10591
rect 16773 10557 16807 10591
rect 18613 10557 18647 10591
rect 19625 10557 19659 10591
rect 22569 10557 22603 10591
rect 25605 10557 25639 10591
rect 10149 10489 10183 10523
rect 15669 10489 15703 10523
rect 21189 10489 21223 10523
rect 21925 10489 21959 10523
rect 22937 10489 22971 10523
rect 25053 10489 25087 10523
rect 30757 10489 30791 10523
rect 8217 10421 8251 10455
rect 9045 10421 9079 10455
rect 17601 10421 17635 10455
rect 18981 10421 19015 10455
rect 19533 10421 19567 10455
rect 20453 10421 20487 10455
rect 24041 10421 24075 10455
rect 27169 10421 27203 10455
rect 31401 10421 31435 10455
rect 6653 10217 6687 10251
rect 7941 10217 7975 10251
rect 10011 10217 10045 10251
rect 11529 10217 11563 10251
rect 17509 10217 17543 10251
rect 18705 10217 18739 10251
rect 19422 10217 19456 10251
rect 19717 10217 19751 10251
rect 23857 10217 23891 10251
rect 26249 10217 26283 10251
rect 14473 10149 14507 10183
rect 16865 10149 16899 10183
rect 19533 10149 19567 10183
rect 28825 10149 28859 10183
rect 6009 10081 6043 10115
rect 7573 10081 7607 10115
rect 14105 10081 14139 10115
rect 15577 10081 15611 10115
rect 18337 10081 18371 10115
rect 19625 10081 19659 10115
rect 21465 10081 21499 10115
rect 26985 10081 27019 10115
rect 5181 10013 5215 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6561 10013 6595 10047
rect 7757 10013 7791 10047
rect 9137 10013 9171 10047
rect 9781 10013 9815 10047
rect 10977 10013 11011 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 12173 10013 12207 10047
rect 12449 10013 12483 10047
rect 14289 10013 14323 10047
rect 15301 10013 15335 10047
rect 18521 10013 18555 10047
rect 21189 10013 21223 10047
rect 22477 10013 22511 10047
rect 24869 10013 24903 10047
rect 26709 10013 26743 10047
rect 27997 10013 28031 10047
rect 29009 10013 29043 10047
rect 29561 10013 29595 10047
rect 29745 10013 29779 10047
rect 30389 10013 30423 10047
rect 31033 10013 31067 10047
rect 31677 10013 31711 10047
rect 9321 9945 9355 9979
rect 11253 9945 11287 9979
rect 16681 9945 16715 9979
rect 17417 9945 17451 9979
rect 19257 9945 19291 9979
rect 20545 9945 20579 9979
rect 20729 9945 20763 9979
rect 22722 9945 22756 9979
rect 25136 9945 25170 9979
rect 28181 9945 28215 9979
rect 28365 9945 28399 9979
rect 4997 9877 5031 9911
rect 7021 9877 7055 9911
rect 11897 9877 11931 9911
rect 29653 9877 29687 9911
rect 30205 9877 30239 9911
rect 30849 9877 30883 9911
rect 31493 9877 31527 9911
rect 8217 9673 8251 9707
rect 21005 9673 21039 9707
rect 27997 9673 28031 9707
rect 30021 9673 30055 9707
rect 7941 9605 7975 9639
rect 10793 9605 10827 9639
rect 11805 9605 11839 9639
rect 12521 9605 12555 9639
rect 18429 9605 18463 9639
rect 21833 9605 21867 9639
rect 22753 9605 22787 9639
rect 22969 9605 23003 9639
rect 25329 9605 25363 9639
rect 26065 9605 26099 9639
rect 26281 9605 26315 9639
rect 27169 9605 27203 9639
rect 27261 9605 27295 9639
rect 3893 9537 3927 9571
rect 4353 9537 4387 9571
rect 4620 9537 4654 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6929 9537 6963 9571
rect 7665 9537 7699 9571
rect 7849 9537 7883 9571
rect 8079 9537 8113 9571
rect 8769 9537 8803 9571
rect 11621 9537 11655 9571
rect 14473 9537 14507 9571
rect 15577 9537 15611 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 17693 9537 17727 9571
rect 18153 9537 18187 9571
rect 18337 9537 18371 9571
rect 18521 9537 18555 9571
rect 19881 9537 19915 9571
rect 22017 9537 22051 9571
rect 24968 9537 25002 9571
rect 25054 9537 25088 9571
rect 25237 9537 25271 9571
rect 25426 9537 25460 9571
rect 26985 9537 27019 9571
rect 27353 9537 27387 9571
rect 28181 9537 28215 9571
rect 28908 9537 28942 9571
rect 30481 9537 30515 9571
rect 30665 9537 30699 9571
rect 31309 9537 31343 9571
rect 32321 9537 32355 9571
rect 32965 9537 32999 9571
rect 33609 9537 33643 9571
rect 6837 9469 6871 9503
rect 8953 9469 8987 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 12265 9469 12299 9503
rect 14565 9469 14599 9503
rect 15301 9469 15335 9503
rect 19625 9469 19659 9503
rect 22293 9469 22327 9503
rect 23581 9469 23615 9503
rect 23857 9469 23891 9503
rect 28641 9469 28675 9503
rect 10977 9401 11011 9435
rect 14841 9401 14875 9435
rect 23121 9401 23155 9435
rect 26433 9401 26467 9435
rect 3709 9333 3743 9367
rect 5733 9333 5767 9367
rect 13645 9333 13679 9367
rect 14657 9333 14691 9367
rect 17509 9333 17543 9367
rect 18705 9333 18739 9367
rect 22201 9333 22235 9367
rect 22937 9333 22971 9367
rect 25605 9333 25639 9367
rect 26249 9333 26283 9367
rect 27537 9333 27571 9367
rect 30481 9333 30515 9367
rect 31125 9333 31159 9367
rect 32137 9333 32171 9367
rect 32781 9333 32815 9367
rect 33425 9333 33459 9367
rect 7021 9129 7055 9163
rect 13553 9129 13587 9163
rect 18705 9129 18739 9163
rect 19349 9129 19383 9163
rect 19993 9129 20027 9163
rect 25881 9129 25915 9163
rect 28181 9129 28215 9163
rect 30849 9129 30883 9163
rect 17693 9061 17727 9095
rect 33425 9061 33459 9095
rect 9321 8993 9355 9027
rect 14289 8993 14323 9027
rect 24501 8993 24535 9027
rect 28917 8993 28951 9027
rect 2513 8925 2547 8959
rect 4077 8925 4111 8959
rect 6469 8925 6503 8959
rect 6837 8925 6871 8959
rect 7665 8925 7699 8959
rect 8401 8925 8435 8959
rect 9045 8925 9079 8959
rect 9137 8925 9171 8959
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 11759 8925 11793 8959
rect 12541 8925 12575 8959
rect 13001 8925 13035 8959
rect 13277 8925 13311 8959
rect 13369 8925 13403 8959
rect 16313 8925 16347 8959
rect 18153 8925 18187 8959
rect 18429 8925 18463 8959
rect 18521 8925 18555 8959
rect 19533 8925 19567 8959
rect 19993 8925 20027 8959
rect 20177 8925 20211 8959
rect 20269 8925 20303 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 22293 8925 22327 8959
rect 22569 8925 22603 8959
rect 23673 8925 23707 8959
rect 24768 8925 24802 8959
rect 26801 8925 26835 8959
rect 26985 8925 27019 8959
rect 27169 8925 27203 8959
rect 27813 8925 27847 8959
rect 28733 8925 28767 8959
rect 29561 8925 29595 8959
rect 29745 8925 29779 8959
rect 30389 8925 30423 8959
rect 31033 8925 31067 8959
rect 31493 8925 31527 8959
rect 31677 8925 31711 8959
rect 32321 8925 32355 8959
rect 32965 8925 32999 8959
rect 33609 8925 33643 8959
rect 4344 8857 4378 8891
rect 6653 8857 6687 8891
rect 6745 8857 6779 8891
rect 8217 8857 8251 8891
rect 11613 8857 11647 8891
rect 13185 8857 13219 8891
rect 14556 8857 14590 8891
rect 16580 8857 16614 8891
rect 18337 8857 18371 8891
rect 21557 8857 21591 8891
rect 21649 8857 21683 8891
rect 22477 8857 22511 8891
rect 27077 8857 27111 8891
rect 27997 8857 28031 8891
rect 31585 8857 31619 8891
rect 2329 8789 2363 8823
rect 5457 8789 5491 8823
rect 7481 8789 7515 8823
rect 11897 8789 11931 8823
rect 12357 8789 12391 8823
rect 15669 8789 15703 8823
rect 20453 8789 20487 8823
rect 22109 8789 22143 8823
rect 23765 8789 23799 8823
rect 27353 8789 27387 8823
rect 29653 8789 29687 8823
rect 30205 8789 30239 8823
rect 32137 8789 32171 8823
rect 32781 8789 32815 8823
rect 1593 8585 1627 8619
rect 3433 8585 3467 8619
rect 4077 8585 4111 8619
rect 5457 8585 5491 8619
rect 6929 8585 6963 8619
rect 10425 8585 10459 8619
rect 14841 8585 14875 8619
rect 19441 8585 19475 8619
rect 25053 8585 25087 8619
rect 29837 8585 29871 8619
rect 30481 8585 30515 8619
rect 34437 8585 34471 8619
rect 6561 8517 6595 8551
rect 10057 8517 10091 8551
rect 11713 8517 11747 8551
rect 12909 8517 12943 8551
rect 17316 8517 17350 8551
rect 19165 8517 19199 8551
rect 21005 8517 21039 8551
rect 24041 8517 24075 8551
rect 24685 8517 24719 8551
rect 24901 8517 24935 8551
rect 30389 8517 30423 8551
rect 1777 8449 1811 8483
rect 2973 8449 3007 8483
rect 3617 8449 3651 8483
rect 4261 8449 4295 8483
rect 4905 8449 4939 8483
rect 5365 8449 5399 8483
rect 5733 8449 5767 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8289 8449 8323 8483
rect 9873 8449 9907 8483
rect 10149 8449 10183 8483
rect 10241 8449 10275 8483
rect 11529 8449 11563 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 12633 8449 12667 8483
rect 12817 8449 12851 8483
rect 13001 8449 13035 8483
rect 13829 8449 13863 8483
rect 14657 8449 14691 8483
rect 15301 8449 15335 8483
rect 17049 8449 17083 8483
rect 18889 8449 18923 8483
rect 19073 8449 19107 8483
rect 19257 8449 19291 8483
rect 20085 8449 20119 8483
rect 20821 8449 20855 8483
rect 20913 8449 20947 8483
rect 21123 8449 21157 8483
rect 22017 8449 22051 8483
rect 23121 8449 23155 8483
rect 25697 8449 25731 8483
rect 26249 8449 26283 8483
rect 26985 8449 27019 8483
rect 27169 8449 27203 8483
rect 27813 8449 27847 8483
rect 27997 8449 28031 8483
rect 28457 8449 28491 8483
rect 28724 8449 28758 8483
rect 31217 8449 31251 8483
rect 32321 8449 32355 8483
rect 33333 8449 33367 8483
rect 33977 8449 34011 8483
rect 34621 8449 34655 8483
rect 35265 8449 35299 8483
rect 5549 8381 5583 8415
rect 13645 8381 13679 8415
rect 14473 8381 14507 8415
rect 15577 8381 15611 8415
rect 21281 8381 21315 8415
rect 23213 8381 23247 8415
rect 23305 8381 23339 8415
rect 27905 8381 27939 8415
rect 2789 8313 2823 8347
rect 4721 8313 4755 8347
rect 7389 8313 7423 8347
rect 19901 8313 19935 8347
rect 24225 8313 24259 8347
rect 25513 8313 25547 8347
rect 27353 8313 27387 8347
rect 31033 8313 31067 8347
rect 32137 8313 32171 8347
rect 33793 8313 33827 8347
rect 35081 8313 35115 8347
rect 5641 8245 5675 8279
rect 9413 8245 9447 8279
rect 12081 8245 12115 8279
rect 13185 8245 13219 8279
rect 14013 8245 14047 8279
rect 18429 8245 18463 8279
rect 20637 8245 20671 8279
rect 21833 8245 21867 8279
rect 22753 8245 22787 8279
rect 24869 8245 24903 8279
rect 26341 8245 26375 8279
rect 33149 8245 33183 8279
rect 5457 8041 5491 8075
rect 14105 8041 14139 8075
rect 16865 8041 16899 8075
rect 18153 8041 18187 8075
rect 19809 8041 19843 8075
rect 21465 8041 21499 8075
rect 23489 8041 23523 8075
rect 26249 8041 26283 8075
rect 33793 8041 33827 8075
rect 25053 7973 25087 8007
rect 32321 7973 32355 8007
rect 5089 7905 5123 7939
rect 8125 7905 8159 7939
rect 14749 7905 14783 7939
rect 16313 7905 16347 7939
rect 27077 7905 27111 7939
rect 30481 7905 30515 7939
rect 1961 7837 1995 7871
rect 2605 7837 2639 7871
rect 3249 7837 3283 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 5273 7837 5307 7871
rect 5917 7837 5951 7871
rect 6193 7837 6227 7871
rect 6285 7837 6319 7871
rect 7297 7837 7331 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 9873 7837 9907 7871
rect 11713 7837 11747 7871
rect 14289 7837 14323 7871
rect 15025 7837 15059 7871
rect 16037 7837 16071 7871
rect 16221 7837 16255 7871
rect 17141 7837 17175 7871
rect 17785 7837 17819 7871
rect 17969 7837 18003 7871
rect 19257 7837 19291 7871
rect 19625 7837 19659 7871
rect 20913 7837 20947 7871
rect 21373 7837 21407 7871
rect 22109 7837 22143 7871
rect 24869 7837 24903 7871
rect 26157 7837 26191 7871
rect 27537 7837 27571 7871
rect 27804 7837 27838 7871
rect 29745 7837 29779 7871
rect 30748 7837 30782 7871
rect 32505 7837 32539 7871
rect 33149 7837 33183 7871
rect 33977 7837 34011 7871
rect 34897 7837 34931 7871
rect 35173 7837 35207 7871
rect 35817 7837 35851 7871
rect 36461 7837 36495 7871
rect 37197 7837 37231 7871
rect 38025 7837 38059 7871
rect 6101 7769 6135 7803
rect 9229 7769 9263 7803
rect 10140 7769 10174 7803
rect 11980 7769 12014 7803
rect 16865 7769 16899 7803
rect 19441 7769 19475 7803
rect 19533 7769 19567 7803
rect 22376 7769 22410 7803
rect 26893 7769 26927 7803
rect 1777 7701 1811 7735
rect 2421 7701 2455 7735
rect 3801 7701 3835 7735
rect 4445 7701 4479 7735
rect 6469 7701 6503 7735
rect 7113 7701 7147 7735
rect 9321 7701 9355 7735
rect 11253 7701 11287 7735
rect 13093 7701 13127 7735
rect 17049 7701 17083 7735
rect 20729 7701 20763 7735
rect 28917 7701 28951 7735
rect 29929 7701 29963 7735
rect 31861 7701 31895 7735
rect 32965 7701 32999 7735
rect 34713 7701 34747 7735
rect 35081 7701 35115 7735
rect 35633 7701 35667 7735
rect 36277 7701 36311 7735
rect 37013 7701 37047 7735
rect 37841 7701 37875 7735
rect 3709 7497 3743 7531
rect 11897 7497 11931 7531
rect 15209 7497 15243 7531
rect 16037 7497 16071 7531
rect 21281 7497 21315 7531
rect 28549 7497 28583 7531
rect 31401 7497 31435 7531
rect 6745 7429 6779 7463
rect 7450 7429 7484 7463
rect 10977 7429 11011 7463
rect 12786 7429 12820 7463
rect 17141 7429 17175 7463
rect 17969 7429 18003 7463
rect 23857 7429 23891 7463
rect 27629 7429 27663 7463
rect 29460 7429 29494 7463
rect 31033 7429 31067 7463
rect 31233 7429 31267 7463
rect 32404 7429 32438 7463
rect 34244 7429 34278 7463
rect 1593 7361 1627 7395
rect 2605 7361 2639 7395
rect 3249 7361 3283 7395
rect 3893 7361 3927 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 10149 7361 10183 7395
rect 10793 7361 10827 7395
rect 11713 7361 11747 7395
rect 14657 7361 14691 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 15025 7361 15059 7395
rect 15853 7361 15887 7395
rect 17785 7361 17819 7395
rect 18153 7361 18187 7395
rect 18797 7361 18831 7395
rect 19441 7361 19475 7395
rect 19901 7361 19935 7395
rect 20168 7361 20202 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 23121 7361 23155 7395
rect 24685 7361 24719 7395
rect 24777 7361 24811 7395
rect 25053 7361 25087 7395
rect 25697 7361 25731 7395
rect 26433 7361 26467 7395
rect 27261 7361 27295 7395
rect 27445 7361 27479 7395
rect 27813 7361 27847 7395
rect 27905 7361 27939 7395
rect 28733 7361 28767 7395
rect 29193 7361 29227 7395
rect 36001 7361 36035 7395
rect 36185 7361 36219 7395
rect 36277 7361 36311 7395
rect 37473 7361 37507 7395
rect 38117 7361 38151 7395
rect 7205 7293 7239 7327
rect 9137 7293 9171 7327
rect 10609 7293 10643 7327
rect 11529 7293 11563 7327
rect 12541 7293 12575 7327
rect 15669 7293 15703 7327
rect 22385 7293 22419 7327
rect 32137 7293 32171 7327
rect 33977 7293 34011 7327
rect 2421 7225 2455 7259
rect 5641 7225 5675 7259
rect 24961 7225 24995 7259
rect 26249 7225 26283 7259
rect 37933 7225 37967 7259
rect 1409 7157 1443 7191
rect 3065 7157 3099 7191
rect 4353 7157 4387 7191
rect 4997 7157 5031 7191
rect 8585 7157 8619 7191
rect 9045 7157 9079 7191
rect 9505 7157 9539 7191
rect 9965 7157 9999 7191
rect 13921 7157 13955 7191
rect 17233 7157 17267 7191
rect 18613 7157 18647 7191
rect 19257 7157 19291 7191
rect 22937 7157 22971 7191
rect 23949 7157 23983 7191
rect 24501 7157 24535 7191
rect 25513 7157 25547 7191
rect 30573 7157 30607 7191
rect 31217 7157 31251 7191
rect 33517 7157 33551 7191
rect 35357 7157 35391 7191
rect 35817 7157 35851 7191
rect 37289 7157 37323 7191
rect 2329 6953 2363 6987
rect 2973 6953 3007 6987
rect 7941 6953 7975 6987
rect 9137 6953 9171 6987
rect 10793 6953 10827 6987
rect 12357 6953 12391 6987
rect 14381 6953 14415 6987
rect 19901 6953 19935 6987
rect 20821 6953 20855 6987
rect 1685 6885 1719 6919
rect 4721 6885 4755 6919
rect 18337 6885 18371 6919
rect 23213 6885 23247 6919
rect 25881 6885 25915 6919
rect 5549 6817 5583 6851
rect 9229 6817 9263 6851
rect 10793 6817 10827 6851
rect 12265 6817 12299 6851
rect 14197 6817 14231 6851
rect 26617 6817 26651 6851
rect 27813 6817 27847 6851
rect 29561 6817 29595 6851
rect 1869 6749 1903 6783
rect 2513 6749 2547 6783
rect 3157 6749 3191 6783
rect 4261 6749 4295 6783
rect 4905 6749 4939 6783
rect 7389 6749 7423 6783
rect 7757 6749 7791 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 10977 6749 11011 6783
rect 12357 6749 12391 6783
rect 13001 6749 13035 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 14381 6749 14415 6783
rect 15025 6749 15059 6783
rect 16957 6749 16991 6783
rect 19533 6749 19567 6783
rect 21557 6749 21591 6783
rect 21741 6749 21775 6783
rect 22385 6749 22419 6783
rect 22569 6749 22603 6783
rect 23029 6749 23063 6783
rect 24501 6749 24535 6783
rect 24768 6749 24802 6783
rect 26801 6749 26835 6783
rect 27005 6727 27039 6761
rect 27537 6749 27571 6783
rect 27721 6749 27755 6783
rect 27910 6749 27944 6783
rect 28549 6749 28583 6783
rect 29828 6749 29862 6783
rect 31953 6749 31987 6783
rect 33885 6749 33919 6783
rect 34069 6749 34103 6783
rect 34713 6749 34747 6783
rect 36737 6749 36771 6783
rect 37013 6749 37047 6783
rect 37657 6749 37691 6783
rect 5794 6681 5828 6715
rect 7573 6681 7607 6715
rect 7665 6681 7699 6715
rect 10701 6681 10735 6715
rect 12081 6681 12115 6715
rect 13185 6681 13219 6715
rect 14105 6681 14139 6715
rect 15292 6681 15326 6715
rect 17202 6681 17236 6715
rect 19717 6681 19751 6715
rect 20729 6681 20763 6715
rect 21833 6681 21867 6715
rect 21925 6681 21959 6715
rect 26617 6681 26651 6715
rect 26893 6681 26927 6715
rect 27813 6681 27847 6715
rect 28733 6681 28767 6715
rect 32220 6681 32254 6715
rect 34980 6681 35014 6715
rect 36553 6681 36587 6715
rect 4077 6613 4111 6647
rect 6929 6613 6963 6647
rect 9597 6613 9631 6647
rect 11161 6613 11195 6647
rect 12541 6613 12575 6647
rect 13553 6613 13587 6647
rect 14565 6613 14599 6647
rect 16405 6613 16439 6647
rect 22569 6613 22603 6647
rect 30941 6613 30975 6647
rect 33333 6613 33367 6647
rect 36093 6613 36127 6647
rect 36921 6613 36955 6647
rect 37473 6613 37507 6647
rect 1685 6409 1719 6443
rect 2973 6409 3007 6443
rect 5641 6409 5675 6443
rect 7205 6409 7239 6443
rect 8401 6409 8435 6443
rect 11713 6409 11747 6443
rect 15485 6409 15519 6443
rect 15945 6409 15979 6443
rect 17049 6409 17083 6443
rect 19441 6409 19475 6443
rect 19993 6409 20027 6443
rect 21189 6409 21223 6443
rect 23765 6409 23799 6443
rect 26249 6409 26283 6443
rect 28365 6409 28399 6443
rect 29653 6409 29687 6443
rect 32781 6409 32815 6443
rect 36553 6409 36587 6443
rect 4528 6341 4562 6375
rect 8033 6341 8067 6375
rect 9312 6341 9346 6375
rect 13001 6341 13035 6375
rect 13185 6341 13219 6375
rect 15117 6341 15151 6375
rect 15209 6341 15243 6375
rect 18328 6341 18362 6375
rect 29285 6341 29319 6375
rect 29485 6341 29519 6375
rect 32413 6341 32447 6375
rect 32613 6341 32647 6375
rect 35440 6341 35474 6375
rect 1869 6273 1903 6307
rect 2513 6273 2547 6307
rect 3157 6273 3191 6307
rect 3801 6273 3835 6307
rect 4261 6273 4295 6307
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 7849 6273 7883 6307
rect 8125 6273 8159 6307
rect 8217 6273 8251 6307
rect 9045 6273 9079 6307
rect 11529 6273 11563 6307
rect 12449 6273 12483 6307
rect 13645 6273 13679 6307
rect 13921 6273 13955 6307
rect 14979 6273 15013 6307
rect 15301 6273 15335 6307
rect 16129 6273 16163 6307
rect 17234 6273 17268 6307
rect 17325 6273 17359 6307
rect 17601 6273 17635 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 22385 6273 22419 6307
rect 22652 6273 22686 6307
rect 24685 6273 24719 6307
rect 25605 6273 25639 6307
rect 26433 6273 26467 6307
rect 27241 6273 27275 6307
rect 30113 6273 30147 6307
rect 30389 6273 30423 6307
rect 31585 6273 31619 6307
rect 37473 6273 37507 6307
rect 38117 6273 38151 6307
rect 6929 6205 6963 6239
rect 13737 6205 13771 6239
rect 18061 6205 18095 6239
rect 24961 6205 24995 6239
rect 25421 6205 25455 6239
rect 26985 6205 27019 6239
rect 33333 6205 33367 6239
rect 33609 6205 33643 6239
rect 35173 6205 35207 6239
rect 2329 6137 2363 6171
rect 20453 6137 20487 6171
rect 3617 6069 3651 6103
rect 6745 6069 6779 6103
rect 10425 6069 10459 6103
rect 12265 6069 12299 6103
rect 13645 6069 13679 6103
rect 14105 6069 14139 6103
rect 17509 6069 17543 6103
rect 24501 6069 24535 6103
rect 24869 6069 24903 6103
rect 25789 6069 25823 6103
rect 29469 6069 29503 6103
rect 31401 6069 31435 6103
rect 32597 6069 32631 6103
rect 37289 6069 37323 6103
rect 37933 6069 37967 6103
rect 1777 5865 1811 5899
rect 5549 5865 5583 5899
rect 12357 5865 12391 5899
rect 15117 5865 15151 5899
rect 18613 5865 18647 5899
rect 21005 5865 21039 5899
rect 23489 5865 23523 5899
rect 25789 5865 25823 5899
rect 27629 5865 27663 5899
rect 29929 5865 29963 5899
rect 32965 5865 32999 5899
rect 33793 5865 33827 5899
rect 33977 5865 34011 5899
rect 35173 5865 35207 5899
rect 35357 5865 35391 5899
rect 2421 5797 2455 5831
rect 8401 5797 8435 5831
rect 13553 5797 13587 5831
rect 17693 5797 17727 5831
rect 22477 5797 22511 5831
rect 30113 5797 30147 5831
rect 33149 5797 33183 5831
rect 4169 5729 4203 5763
rect 10425 5729 10459 5763
rect 15117 5729 15151 5763
rect 19625 5729 19659 5763
rect 23581 5729 23615 5763
rect 31493 5729 31527 5763
rect 31769 5729 31803 5763
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 6377 5661 6411 5695
rect 7481 5661 7515 5695
rect 9321 5661 9355 5695
rect 10977 5661 11011 5695
rect 13369 5661 13403 5695
rect 14381 5661 14415 5695
rect 15301 5661 15335 5695
rect 16221 5661 16255 5695
rect 16497 5661 16531 5695
rect 17417 5661 17451 5695
rect 17509 5661 17543 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 19881 5661 19915 5695
rect 22017 5661 22051 5695
rect 23305 5661 23339 5695
rect 24409 5661 24443 5695
rect 26249 5661 26283 5695
rect 28365 5661 28399 5695
rect 29009 5661 29043 5695
rect 30757 5661 30791 5695
rect 36001 5661 36035 5695
rect 36645 5661 36679 5695
rect 37289 5661 37323 5695
rect 37841 5661 37875 5695
rect 4414 5593 4448 5627
rect 6009 5593 6043 5627
rect 6193 5593 6227 5627
rect 8217 5593 8251 5627
rect 10149 5593 10183 5627
rect 11222 5593 11256 5627
rect 14565 5593 14599 5627
rect 15025 5593 15059 5627
rect 16037 5593 16071 5627
rect 17233 5593 17267 5627
rect 18245 5593 18279 5627
rect 24654 5593 24688 5627
rect 26516 5593 26550 5627
rect 29745 5593 29779 5627
rect 29945 5593 29979 5627
rect 32781 5593 32815 5627
rect 32981 5593 33015 5627
rect 33609 5593 33643 5627
rect 34989 5593 35023 5627
rect 3065 5525 3099 5559
rect 7573 5525 7607 5559
rect 9505 5525 9539 5559
rect 15485 5525 15519 5559
rect 16405 5525 16439 5559
rect 22017 5525 22051 5559
rect 23857 5525 23891 5559
rect 28181 5525 28215 5559
rect 28825 5525 28859 5559
rect 30573 5525 30607 5559
rect 33809 5525 33843 5559
rect 35189 5525 35223 5559
rect 35817 5525 35851 5559
rect 36461 5525 36495 5559
rect 37105 5525 37139 5559
rect 38025 5525 38059 5559
rect 2329 5321 2363 5355
rect 5181 5321 5215 5355
rect 8309 5321 8343 5355
rect 9689 5321 9723 5355
rect 11897 5321 11931 5355
rect 13921 5321 13955 5355
rect 22845 5321 22879 5355
rect 24133 5321 24167 5355
rect 29393 5321 29427 5355
rect 29561 5321 29595 5355
rect 30849 5321 30883 5355
rect 32347 5321 32381 5355
rect 33165 5321 33199 5355
rect 33333 5321 33367 5355
rect 33793 5321 33827 5355
rect 36645 5321 36679 5355
rect 37657 5321 37691 5355
rect 7196 5253 7230 5287
rect 9505 5253 9539 5287
rect 12786 5253 12820 5287
rect 17049 5253 17083 5287
rect 28273 5253 28307 5287
rect 29193 5253 29227 5287
rect 30021 5253 30055 5287
rect 30221 5253 30255 5287
rect 32137 5253 32171 5287
rect 32965 5253 32999 5287
rect 35532 5253 35566 5287
rect 37289 5253 37323 5287
rect 37489 5253 37523 5287
rect 1869 5185 1903 5219
rect 2513 5185 2547 5219
rect 2973 5185 3007 5219
rect 3229 5185 3263 5219
rect 4813 5185 4847 5219
rect 4997 5185 5031 5219
rect 5825 5185 5859 5219
rect 6929 5185 6963 5219
rect 9321 5185 9355 5219
rect 10425 5185 10459 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 12548 5185 12582 5219
rect 15117 5185 15151 5219
rect 15209 5185 15243 5219
rect 15485 5185 15519 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 18981 5185 19015 5219
rect 19717 5185 19751 5219
rect 20729 5185 20763 5219
rect 21833 5185 21867 5219
rect 22017 5185 22051 5219
rect 22201 5185 22235 5219
rect 22661 5185 22695 5219
rect 22937 5185 22971 5219
rect 23397 5185 23431 5219
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 24317 5185 24351 5219
rect 24961 5185 24995 5219
rect 25605 5185 25639 5219
rect 26249 5185 26283 5219
rect 27169 5185 27203 5219
rect 31033 5185 31067 5219
rect 33977 5185 34011 5219
rect 34621 5185 34655 5219
rect 10149 5117 10183 5151
rect 16037 5117 16071 5151
rect 17693 5117 17727 5151
rect 17969 5117 18003 5151
rect 35265 5117 35299 5151
rect 4353 5049 4387 5083
rect 22661 5049 22695 5083
rect 28457 5049 28491 5083
rect 30389 5049 30423 5083
rect 32505 5049 32539 5083
rect 1685 4981 1719 5015
rect 5641 4981 5675 5015
rect 14933 4981 14967 5015
rect 15393 4981 15427 5015
rect 17141 4981 17175 5015
rect 19165 4981 19199 5015
rect 19901 4981 19935 5015
rect 20821 4981 20855 5015
rect 23397 4981 23431 5015
rect 24777 4981 24811 5015
rect 25421 4981 25455 5015
rect 26065 4981 26099 5015
rect 26985 4981 27019 5015
rect 29377 4981 29411 5015
rect 30205 4981 30239 5015
rect 32321 4981 32355 5015
rect 33149 4981 33183 5015
rect 34437 4981 34471 5015
rect 37473 4981 37507 5015
rect 3065 4777 3099 4811
rect 5273 4777 5307 4811
rect 8401 4777 8435 4811
rect 10241 4777 10275 4811
rect 10701 4777 10735 4811
rect 11621 4777 11655 4811
rect 13461 4777 13495 4811
rect 15945 4777 15979 4811
rect 25605 4777 25639 4811
rect 28825 4777 28859 4811
rect 31677 4777 31711 4811
rect 31861 4777 31895 4811
rect 32597 4777 32631 4811
rect 32781 4777 32815 4811
rect 34897 4777 34931 4811
rect 35081 4777 35115 4811
rect 35725 4777 35759 4811
rect 35909 4777 35943 4811
rect 36645 4777 36679 4811
rect 36829 4777 36863 4811
rect 12081 4709 12115 4743
rect 26157 4709 26191 4743
rect 27169 4709 27203 4743
rect 29009 4709 29043 4743
rect 33885 4709 33919 4743
rect 4261 4641 4295 4675
rect 5733 4641 5767 4675
rect 6745 4641 6779 4675
rect 8953 4641 8987 4675
rect 14565 4641 14599 4675
rect 20177 4641 20211 4675
rect 1961 4573 1995 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 3893 4573 3927 4607
rect 5458 4573 5492 4607
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 7021 4573 7055 4607
rect 9229 4573 9263 4607
rect 10408 4573 10442 4607
rect 10518 4573 10552 4607
rect 10793 4573 10827 4607
rect 11805 4573 11839 4607
rect 11897 4573 11931 4607
rect 12173 4573 12207 4607
rect 13185 4573 13219 4607
rect 13337 4573 13371 4607
rect 13553 4573 13587 4607
rect 16405 4573 16439 4607
rect 18521 4573 18555 4607
rect 19809 4573 19843 4607
rect 20637 4573 20671 4607
rect 21373 4573 21407 4607
rect 22109 4573 22143 4607
rect 22845 4573 22879 4607
rect 23581 4573 23615 4607
rect 24593 4573 24627 4607
rect 26341 4573 26375 4607
rect 26893 4573 26927 4607
rect 26985 4573 27019 4607
rect 27813 4573 27847 4607
rect 29561 4573 29595 4607
rect 29745 4573 29779 4607
rect 30021 4573 30055 4607
rect 30757 4573 30791 4607
rect 31033 4573 31067 4607
rect 33425 4573 33459 4607
rect 34069 4573 34103 4607
rect 37841 4573 37875 4607
rect 28871 4539 28905 4573
rect 4077 4505 4111 4539
rect 8033 4505 8067 4539
rect 8217 4505 8251 4539
rect 14810 4505 14844 4539
rect 16589 4505 16623 4539
rect 16773 4505 16807 4539
rect 17325 4505 17359 4539
rect 17509 4505 17543 4539
rect 18153 4505 18187 4539
rect 18337 4505 18371 4539
rect 19993 4505 20027 4539
rect 25513 4505 25547 4539
rect 28641 4505 28675 4539
rect 30941 4505 30975 4539
rect 31493 4505 31527 4539
rect 32413 4505 32447 4539
rect 32629 4505 32663 4539
rect 34713 4505 34747 4539
rect 34913 4505 34947 4539
rect 35541 4505 35575 4539
rect 36461 4505 36495 4539
rect 36661 4505 36695 4539
rect 1777 4437 1811 4471
rect 2421 4437 2455 4471
rect 13001 4437 13035 4471
rect 17693 4437 17727 4471
rect 20821 4437 20855 4471
rect 21557 4437 21591 4471
rect 22293 4437 22327 4471
rect 23029 4437 23063 4471
rect 23765 4437 23799 4471
rect 24409 4437 24443 4471
rect 27629 4437 27663 4471
rect 29929 4437 29963 4471
rect 30573 4437 30607 4471
rect 31703 4437 31737 4471
rect 33241 4437 33275 4471
rect 35741 4437 35775 4471
rect 38025 4437 38059 4471
rect 2881 4233 2915 4267
rect 3525 4233 3559 4267
rect 7481 4233 7515 4267
rect 11897 4233 11931 4267
rect 13645 4233 13679 4267
rect 20453 4233 20487 4267
rect 27353 4233 27387 4267
rect 29561 4233 29595 4267
rect 35557 4233 35591 4267
rect 11529 4165 11563 4199
rect 12817 4165 12851 4199
rect 13001 4165 13035 4199
rect 35357 4165 35391 4199
rect 1869 4097 1903 4131
rect 3065 4097 3099 4131
rect 3709 4097 3743 4131
rect 4169 4097 4203 4131
rect 4353 4097 4387 4131
rect 4445 4097 4479 4131
rect 4721 4097 4755 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 5549 4097 5583 4131
rect 5825 4097 5859 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 6929 4097 6963 4131
rect 7665 4097 7699 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 11713 4097 11747 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 14473 4097 14507 4131
rect 14565 4097 14599 4131
rect 14841 4097 14875 4131
rect 16865 4097 16899 4131
rect 17325 4097 17359 4131
rect 18880 4097 18914 4131
rect 20637 4097 20671 4131
rect 20729 4097 20763 4131
rect 21005 4097 21039 4131
rect 22293 4097 22327 4131
rect 22560 4097 22594 4131
rect 24409 4097 24443 4131
rect 24593 4097 24627 4131
rect 25053 4097 25087 4131
rect 25237 4097 25271 4131
rect 25421 4097 25455 4131
rect 26249 4097 26283 4131
rect 26433 4097 26467 4131
rect 26985 4097 27019 4131
rect 27169 4097 27203 4131
rect 28181 4097 28215 4131
rect 28448 4097 28482 4131
rect 30021 4097 30055 4131
rect 30288 4097 30322 4131
rect 32321 4097 32355 4131
rect 32505 4097 32539 4131
rect 32597 4097 32631 4131
rect 33784 4097 33818 4131
rect 36461 4097 36495 4131
rect 37289 4097 37323 4131
rect 4629 4029 4663 4063
rect 8493 4029 8527 4063
rect 9781 4029 9815 4063
rect 10057 4029 10091 4063
rect 14749 4029 14783 4063
rect 15301 4029 15335 4063
rect 15577 4029 15611 4063
rect 17601 4029 17635 4063
rect 18613 4029 18647 4063
rect 20913 4029 20947 4063
rect 24225 4029 24259 4063
rect 26065 4029 26099 4063
rect 33517 4029 33551 4063
rect 35725 3961 35759 3995
rect 36645 3961 36679 3995
rect 1685 3893 1719 3927
rect 5733 3893 5767 3927
rect 6377 3893 6411 3927
rect 6837 3893 6871 3927
rect 7941 3893 7975 3927
rect 8723 3893 8757 3927
rect 14289 3893 14323 3927
rect 16681 3893 16715 3927
rect 19993 3893 20027 3927
rect 23673 3893 23707 3927
rect 31401 3893 31435 3927
rect 32137 3893 32171 3927
rect 34897 3893 34931 3927
rect 35541 3893 35575 3927
rect 37473 3893 37507 3927
rect 7021 3689 7055 3723
rect 17233 3689 17267 3723
rect 17877 3689 17911 3723
rect 19257 3689 19291 3723
rect 20361 3689 20395 3723
rect 25697 3689 25731 3723
rect 27905 3689 27939 3723
rect 32413 3689 32447 3723
rect 33977 3689 34011 3723
rect 34161 3689 34195 3723
rect 36093 3689 36127 3723
rect 36737 3689 36771 3723
rect 36921 3689 36955 3723
rect 2329 3621 2363 3655
rect 5181 3621 5215 3655
rect 8033 3621 8067 3655
rect 10333 3621 10367 3655
rect 12357 3621 12391 3655
rect 17601 3621 17635 3655
rect 25605 3621 25639 3655
rect 26525 3621 26559 3655
rect 27813 3621 27847 3655
rect 37565 3621 37599 3655
rect 14565 3553 14599 3587
rect 15853 3553 15887 3587
rect 18337 3553 18371 3587
rect 20913 3553 20947 3587
rect 24777 3553 24811 3587
rect 26157 3553 26191 3587
rect 27445 3553 27479 3587
rect 29837 3553 29871 3587
rect 31033 3553 31067 3587
rect 34713 3553 34747 3587
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 1961 3485 1995 3519
rect 3249 3485 3283 3519
rect 3801 3485 3835 3519
rect 5641 3485 5675 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 8125 3485 8159 3519
rect 8953 3485 8987 3519
rect 10977 3485 11011 3519
rect 11244 3485 11278 3519
rect 13001 3485 13035 3519
rect 14272 3485 14306 3519
rect 14381 3485 14415 3519
rect 14657 3485 14691 3519
rect 16109 3485 16143 3519
rect 18061 3485 18095 3519
rect 18153 3485 18187 3519
rect 18429 3485 18463 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20177 3485 20211 3519
rect 20453 3485 20487 3519
rect 22845 3485 22879 3519
rect 23029 3485 23063 3519
rect 23213 3485 23247 3519
rect 23857 3485 23891 3519
rect 24409 3485 24443 3519
rect 24593 3485 24627 3519
rect 28641 3485 28675 3519
rect 28917 3485 28951 3519
rect 29561 3485 29595 3519
rect 33057 3485 33091 3519
rect 33333 3485 33367 3519
rect 37381 3485 37415 3519
rect 34023 3451 34057 3485
rect 4046 3417 4080 3451
rect 5886 3417 5920 3451
rect 7573 3417 7607 3451
rect 9198 3417 9232 3451
rect 12817 3417 12851 3451
rect 13185 3417 13219 3451
rect 15117 3417 15151 3451
rect 15301 3417 15335 3451
rect 21180 3417 21214 3451
rect 25237 3417 25271 3451
rect 31300 3417 31334 3451
rect 33241 3417 33275 3451
rect 33793 3417 33827 3451
rect 34980 3417 35014 3451
rect 36553 3417 36587 3451
rect 3065 3349 3099 3383
rect 14105 3349 14139 3383
rect 15485 3349 15519 3383
rect 19901 3349 19935 3383
rect 22293 3349 22327 3383
rect 23673 3349 23707 3383
rect 26617 3349 26651 3383
rect 28457 3349 28491 3383
rect 28825 3349 28859 3383
rect 32873 3349 32907 3383
rect 36753 3349 36787 3383
rect 2329 3145 2363 3179
rect 2973 3145 3007 3179
rect 3985 3145 4019 3179
rect 8125 3145 8159 3179
rect 15761 3145 15795 3179
rect 23029 3145 23063 3179
rect 23857 3145 23891 3179
rect 25329 3145 25363 3179
rect 26157 3145 26191 3179
rect 29101 3145 29135 3179
rect 31309 3145 31343 3179
rect 33517 3145 33551 3179
rect 35005 3145 35039 3179
rect 35173 3145 35207 3179
rect 36185 3145 36219 3179
rect 3617 3077 3651 3111
rect 3801 3077 3835 3111
rect 5457 3077 5491 3111
rect 7001 3077 7035 3111
rect 29561 3077 29595 3111
rect 29761 3077 29795 3111
rect 32404 3077 32438 3111
rect 34805 3077 34839 3111
rect 35817 3077 35851 3111
rect 36017 3077 36051 3111
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 3157 3009 3191 3043
rect 4629 3009 4663 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5641 3009 5675 3043
rect 6745 3009 6779 3043
rect 8769 3009 8803 3043
rect 8861 3009 8895 3043
rect 9137 3009 9171 3043
rect 9597 3009 9631 3043
rect 9853 3009 9887 3043
rect 11713 3009 11747 3043
rect 11805 3009 11839 3043
rect 12081 3009 12115 3043
rect 12541 3009 12575 3043
rect 12797 3009 12831 3043
rect 14381 3009 14415 3043
rect 14637 3009 14671 3043
rect 17049 3009 17083 3043
rect 17305 3009 17339 3043
rect 19073 3009 19107 3043
rect 19165 3009 19199 3043
rect 19395 3009 19429 3043
rect 19901 3009 19935 3043
rect 20168 3009 20202 3043
rect 22017 3009 22051 3043
rect 22753 3009 22787 3043
rect 22845 3009 22879 3043
rect 23673 3009 23707 3043
rect 24501 3009 24535 3043
rect 24961 3009 24995 3043
rect 25145 3009 25179 3043
rect 25973 3009 26007 3043
rect 26985 3009 27019 3043
rect 27721 3009 27755 3043
rect 27988 3009 28022 3043
rect 30389 3009 30423 3043
rect 31125 3009 31159 3043
rect 32137 3009 32171 3043
rect 33977 3009 34011 3043
rect 37289 3009 37323 3043
rect 11529 2941 11563 2975
rect 21833 2941 21867 2975
rect 23489 2941 23523 2975
rect 25789 2941 25823 2975
rect 4445 2873 4479 2907
rect 10977 2873 11011 2907
rect 11989 2873 12023 2907
rect 13921 2873 13955 2907
rect 18429 2873 18463 2907
rect 22201 2873 22235 2907
rect 27169 2873 27203 2907
rect 29929 2873 29963 2907
rect 37473 2873 37507 2907
rect 1685 2805 1719 2839
rect 4905 2805 4939 2839
rect 5825 2805 5859 2839
rect 8585 2805 8619 2839
rect 9045 2805 9079 2839
rect 18889 2805 18923 2839
rect 19349 2805 19383 2839
rect 21281 2805 21315 2839
rect 24317 2805 24351 2839
rect 29745 2805 29779 2839
rect 30573 2805 30607 2839
rect 34161 2805 34195 2839
rect 34989 2805 35023 2839
rect 36001 2805 36035 2839
rect 5641 2601 5675 2635
rect 6745 2601 6779 2635
rect 8217 2601 8251 2635
rect 9965 2601 9999 2635
rect 11621 2601 11655 2635
rect 14473 2601 14507 2635
rect 18061 2601 18095 2635
rect 19625 2601 19659 2635
rect 20545 2601 20579 2635
rect 30481 2601 30515 2635
rect 33793 2601 33827 2635
rect 4997 2533 5031 2567
rect 15301 2533 15335 2567
rect 17325 2533 17359 2567
rect 18521 2533 18555 2567
rect 25789 2533 25823 2567
rect 32321 2533 32355 2567
rect 34897 2533 34931 2567
rect 36369 2533 36403 2567
rect 3249 2465 3283 2499
rect 7757 2465 7791 2499
rect 9321 2465 9355 2499
rect 10425 2465 10459 2499
rect 24777 2465 24811 2499
rect 25145 2465 25179 2499
rect 27261 2465 27295 2499
rect 3801 2397 3835 2431
rect 5181 2397 5215 2431
rect 5825 2397 5859 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 8401 2397 8435 2431
rect 8953 2397 8987 2431
rect 10149 2397 10183 2431
rect 10241 2397 10275 2431
rect 10517 2397 10551 2431
rect 11805 2397 11839 2431
rect 12449 2397 12483 2431
rect 13093 2397 13127 2431
rect 14657 2397 14691 2431
rect 15117 2397 15151 2431
rect 15853 2397 15887 2431
rect 17141 2397 17175 2431
rect 18245 2397 18279 2431
rect 18337 2397 18371 2431
rect 18613 2397 18647 2431
rect 19257 2397 19291 2431
rect 19441 2397 19475 2431
rect 20177 2397 20211 2431
rect 21005 2397 21039 2431
rect 22109 2397 22143 2431
rect 22385 2397 22419 2431
rect 23581 2397 23615 2431
rect 24961 2397 24995 2431
rect 25605 2397 25639 2431
rect 26985 2397 27019 2431
rect 28273 2397 28307 2431
rect 29561 2397 29595 2431
rect 30297 2397 30331 2431
rect 31033 2397 31067 2431
rect 32137 2397 32171 2431
rect 32873 2397 32907 2431
rect 33609 2397 33643 2431
rect 34713 2397 34747 2431
rect 35449 2397 35483 2431
rect 36185 2397 36219 2431
rect 1869 2329 1903 2363
rect 2053 2329 2087 2363
rect 7573 2329 7607 2363
rect 9137 2329 9171 2363
rect 12909 2329 12943 2363
rect 20361 2329 20395 2363
rect 37933 2329 37967 2363
rect 3985 2261 4019 2295
rect 12265 2261 12299 2295
rect 13277 2261 13311 2295
rect 16037 2261 16071 2295
rect 21189 2261 21223 2295
rect 23765 2261 23799 2295
rect 28457 2261 28491 2295
rect 29745 2261 29779 2295
rect 31217 2261 31251 2295
rect 33057 2261 33091 2295
rect 35633 2261 35667 2295
rect 38025 2261 38059 2295
<< metal1 >>
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 15194 47240 15200 47252
rect 15155 47212 15200 47240
rect 15194 47200 15200 47212
rect 15252 47200 15258 47252
rect 25222 47240 25228 47252
rect 25183 47212 25228 47240
rect 25222 47200 25228 47212
rect 25280 47200 25286 47252
rect 35253 47243 35311 47249
rect 35253 47209 35265 47243
rect 35299 47240 35311 47243
rect 35342 47240 35348 47252
rect 35299 47212 35348 47240
rect 35299 47209 35311 47212
rect 35253 47203 35311 47209
rect 35342 47200 35348 47212
rect 35400 47200 35406 47252
rect 5074 47036 5080 47048
rect 5035 47008 5080 47036
rect 5074 46996 5080 47008
rect 5132 46996 5138 47048
rect 15013 47039 15071 47045
rect 15013 47005 15025 47039
rect 15059 47036 15071 47039
rect 19242 47036 19248 47048
rect 15059 47008 19248 47036
rect 15059 47005 15071 47008
rect 15013 46999 15071 47005
rect 19242 46996 19248 47008
rect 19300 46996 19306 47048
rect 24854 46996 24860 47048
rect 24912 47036 24918 47048
rect 25041 47039 25099 47045
rect 25041 47036 25053 47039
rect 24912 47008 25053 47036
rect 24912 46996 24918 47008
rect 25041 47005 25053 47008
rect 25087 47005 25099 47039
rect 25041 46999 25099 47005
rect 35069 47039 35127 47045
rect 35069 47005 35081 47039
rect 35115 47036 35127 47039
rect 35342 47036 35348 47048
rect 35115 47008 35348 47036
rect 35115 47005 35127 47008
rect 35069 46999 35127 47005
rect 35342 46996 35348 47008
rect 35400 46996 35406 47048
rect 5258 46900 5264 46912
rect 5219 46872 5264 46900
rect 5258 46860 5264 46872
rect 5316 46860 5322 46912
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 19242 46656 19248 46708
rect 19300 46696 19306 46708
rect 19797 46699 19855 46705
rect 19797 46696 19809 46699
rect 19300 46668 19809 46696
rect 19300 46656 19306 46668
rect 19797 46665 19809 46668
rect 19843 46665 19855 46699
rect 19797 46659 19855 46665
rect 19981 46563 20039 46569
rect 19981 46529 19993 46563
rect 20027 46560 20039 46563
rect 20530 46560 20536 46572
rect 20027 46532 20536 46560
rect 20027 46529 20039 46532
rect 19981 46523 20039 46529
rect 20530 46520 20536 46532
rect 20588 46520 20594 46572
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30716 19487 30719
rect 20990 30716 20996 30728
rect 19475 30688 20996 30716
rect 19475 30685 19487 30688
rect 19429 30679 19487 30685
rect 20990 30676 20996 30688
rect 21048 30676 21054 30728
rect 19242 30580 19248 30592
rect 19203 30552 19248 30580
rect 19242 30540 19248 30552
rect 19300 30540 19306 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 19242 30317 19248 30320
rect 19236 30308 19248 30317
rect 17144 30280 19012 30308
rect 19203 30280 19248 30308
rect 15746 30200 15752 30252
rect 15804 30240 15810 30252
rect 17144 30249 17172 30280
rect 17129 30243 17187 30249
rect 17129 30240 17141 30243
rect 15804 30212 17141 30240
rect 15804 30200 15810 30212
rect 17129 30209 17141 30212
rect 17175 30209 17187 30243
rect 17129 30203 17187 30209
rect 17396 30243 17454 30249
rect 17396 30209 17408 30243
rect 17442 30240 17454 30243
rect 18414 30240 18420 30252
rect 17442 30212 18420 30240
rect 17442 30209 17454 30212
rect 17396 30203 17454 30209
rect 18414 30200 18420 30212
rect 18472 30200 18478 30252
rect 18984 30249 19012 30280
rect 19236 30271 19248 30280
rect 19242 30268 19248 30271
rect 19300 30268 19306 30320
rect 18969 30243 19027 30249
rect 18969 30209 18981 30243
rect 19015 30209 19027 30243
rect 18969 30203 19027 30209
rect 18506 30036 18512 30048
rect 18467 30008 18512 30036
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 20349 30039 20407 30045
rect 20349 30005 20361 30039
rect 20395 30036 20407 30039
rect 20438 30036 20444 30048
rect 20395 30008 20444 30036
rect 20395 30005 20407 30008
rect 20349 29999 20407 30005
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 18414 29832 18420 29844
rect 18375 29804 18420 29832
rect 18414 29792 18420 29804
rect 18472 29792 18478 29844
rect 20990 29832 20996 29844
rect 20951 29804 20996 29832
rect 20990 29792 20996 29804
rect 21048 29792 21054 29844
rect 15746 29696 15752 29708
rect 15707 29668 15752 29696
rect 15746 29656 15752 29668
rect 15804 29656 15810 29708
rect 19797 29699 19855 29705
rect 19797 29696 19809 29699
rect 17604 29668 19809 29696
rect 17604 29640 17632 29668
rect 19797 29665 19809 29668
rect 19843 29696 19855 29699
rect 20622 29696 20628 29708
rect 19843 29668 20628 29696
rect 19843 29665 19855 29668
rect 19797 29659 19855 29665
rect 20622 29656 20628 29668
rect 20680 29656 20686 29708
rect 17586 29628 17592 29640
rect 17547 29600 17592 29628
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 17770 29628 17776 29640
rect 17731 29600 17776 29628
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18601 29631 18659 29637
rect 18601 29628 18613 29631
rect 18003 29600 18613 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 18601 29597 18613 29600
rect 18647 29597 18659 29631
rect 19978 29628 19984 29640
rect 19939 29600 19984 29628
rect 18601 29591 18659 29597
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 20806 29628 20812 29640
rect 20767 29600 20812 29628
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 16016 29563 16074 29569
rect 16016 29529 16028 29563
rect 16062 29560 16074 29563
rect 16666 29560 16672 29572
rect 16062 29532 16672 29560
rect 16062 29529 16074 29532
rect 16016 29523 16074 29529
rect 16666 29520 16672 29532
rect 16724 29520 16730 29572
rect 17129 29495 17187 29501
rect 17129 29461 17141 29495
rect 17175 29492 17187 29495
rect 17402 29492 17408 29504
rect 17175 29464 17408 29492
rect 17175 29461 17187 29464
rect 17129 29455 17187 29461
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 20165 29495 20223 29501
rect 20165 29461 20177 29495
rect 20211 29492 20223 29495
rect 21266 29492 21272 29504
rect 20211 29464 21272 29492
rect 20211 29461 20223 29464
rect 20165 29455 20223 29461
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 16666 29288 16672 29300
rect 16627 29260 16672 29288
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 17770 29248 17776 29300
rect 17828 29288 17834 29300
rect 18417 29291 18475 29297
rect 18417 29288 18429 29291
rect 17828 29260 18429 29288
rect 17828 29248 17834 29260
rect 18417 29257 18429 29260
rect 18463 29257 18475 29291
rect 18417 29251 18475 29257
rect 19429 29291 19487 29297
rect 19429 29257 19441 29291
rect 19475 29288 19487 29291
rect 20806 29288 20812 29300
rect 19475 29260 20812 29288
rect 19475 29257 19487 29260
rect 19429 29251 19487 29257
rect 20806 29248 20812 29260
rect 20864 29248 20870 29300
rect 21821 29291 21879 29297
rect 21821 29257 21833 29291
rect 21867 29257 21879 29291
rect 21821 29251 21879 29257
rect 19153 29223 19211 29229
rect 17880 29192 18920 29220
rect 15930 29152 15936 29164
rect 15891 29124 15936 29152
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 17880 29161 17908 29192
rect 17865 29155 17923 29161
rect 17865 29121 17877 29155
rect 17911 29121 17923 29155
rect 18046 29152 18052 29164
rect 18007 29124 18052 29152
rect 17865 29115 17923 29121
rect 17880 29084 17908 29115
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 18892 29161 18920 29192
rect 19153 29189 19165 29223
rect 19199 29220 19211 29223
rect 20156 29223 20214 29229
rect 19199 29192 19840 29220
rect 19199 29189 19211 29192
rect 19153 29183 19211 29189
rect 18141 29155 18199 29161
rect 18141 29121 18153 29155
rect 18187 29121 18199 29155
rect 18141 29115 18199 29121
rect 18279 29155 18337 29161
rect 18279 29121 18291 29155
rect 18325 29152 18337 29155
rect 18877 29155 18935 29161
rect 18325 29124 18460 29152
rect 18325 29121 18337 29124
rect 18279 29115 18337 29121
rect 17954 29084 17960 29096
rect 17880 29056 17960 29084
rect 17954 29044 17960 29056
rect 18012 29044 18018 29096
rect 18156 29016 18184 29115
rect 18432 29096 18460 29124
rect 18877 29121 18889 29155
rect 18923 29121 18935 29155
rect 19058 29152 19064 29164
rect 19019 29124 19064 29152
rect 18877 29115 18935 29121
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 19242 29152 19248 29164
rect 19168 29124 19248 29152
rect 18414 29044 18420 29096
rect 18472 29084 18478 29096
rect 19168 29084 19196 29124
rect 19242 29112 19248 29124
rect 19300 29112 19306 29164
rect 19812 29152 19840 29192
rect 20156 29189 20168 29223
rect 20202 29220 20214 29223
rect 21836 29220 21864 29251
rect 20202 29192 21864 29220
rect 20202 29189 20214 29192
rect 20156 29183 20214 29189
rect 20438 29152 20444 29164
rect 19812 29124 20444 29152
rect 20438 29112 20444 29124
rect 20496 29112 20502 29164
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22646 29152 22652 29164
rect 22051 29124 22652 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 19886 29084 19892 29096
rect 18472 29056 19196 29084
rect 19847 29056 19892 29084
rect 18472 29044 18478 29056
rect 19886 29044 19892 29056
rect 19944 29044 19950 29096
rect 18506 29016 18512 29028
rect 18156 28988 18512 29016
rect 18506 28976 18512 28988
rect 18564 29016 18570 29028
rect 19150 29016 19156 29028
rect 18564 28988 19156 29016
rect 18564 28976 18570 28988
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 21269 29019 21327 29025
rect 21269 28985 21281 29019
rect 21315 28985 21327 29019
rect 21269 28979 21327 28985
rect 15749 28951 15807 28957
rect 15749 28917 15761 28951
rect 15795 28948 15807 28951
rect 16114 28948 16120 28960
rect 15795 28920 16120 28948
rect 15795 28917 15807 28920
rect 15749 28911 15807 28917
rect 16114 28908 16120 28920
rect 16172 28908 16178 28960
rect 20806 28908 20812 28960
rect 20864 28948 20870 28960
rect 21284 28948 21312 28979
rect 20864 28920 21312 28948
rect 20864 28908 20870 28920
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 19797 28747 19855 28753
rect 19797 28713 19809 28747
rect 19843 28744 19855 28747
rect 19978 28744 19984 28756
rect 19843 28716 19984 28744
rect 19843 28713 19855 28716
rect 19797 28707 19855 28713
rect 19978 28704 19984 28716
rect 20036 28704 20042 28756
rect 20622 28704 20628 28756
rect 20680 28744 20686 28756
rect 22646 28744 22652 28756
rect 20680 28716 22094 28744
rect 22607 28716 22652 28744
rect 20680 28704 20686 28716
rect 15746 28568 15752 28620
rect 15804 28608 15810 28620
rect 15841 28611 15899 28617
rect 15841 28608 15853 28611
rect 15804 28580 15853 28608
rect 15804 28568 15810 28580
rect 15841 28577 15853 28580
rect 15887 28577 15899 28611
rect 17954 28608 17960 28620
rect 15841 28571 15899 28577
rect 17696 28580 17960 28608
rect 16114 28549 16120 28552
rect 16108 28540 16120 28549
rect 16075 28512 16120 28540
rect 16108 28503 16120 28512
rect 16114 28500 16120 28503
rect 16172 28500 16178 28552
rect 17696 28549 17724 28580
rect 17954 28568 17960 28580
rect 18012 28608 18018 28620
rect 22066 28608 22094 28716
rect 22646 28704 22652 28716
rect 22704 28704 22710 28756
rect 22281 28611 22339 28617
rect 22281 28608 22293 28611
rect 18012 28580 19288 28608
rect 22066 28580 22293 28608
rect 18012 28568 18018 28580
rect 17681 28543 17739 28549
rect 17681 28509 17693 28543
rect 17727 28509 17739 28543
rect 17681 28503 17739 28509
rect 18049 28543 18107 28549
rect 18049 28509 18061 28543
rect 18095 28540 18107 28543
rect 18138 28540 18144 28552
rect 18095 28512 18144 28540
rect 18095 28509 18107 28512
rect 18049 28503 18107 28509
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 19260 28549 19288 28580
rect 22281 28577 22293 28580
rect 22327 28577 22339 28611
rect 22281 28571 22339 28577
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19613 28543 19671 28549
rect 19613 28540 19625 28543
rect 19392 28512 19625 28540
rect 19392 28500 19398 28512
rect 19613 28509 19625 28512
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 19944 28512 20453 28540
rect 19944 28500 19950 28512
rect 20441 28509 20453 28512
rect 20487 28540 20499 28543
rect 22094 28540 22100 28552
rect 20487 28512 22100 28540
rect 20487 28509 20499 28512
rect 20441 28503 20499 28509
rect 22094 28500 22100 28512
rect 22152 28500 22158 28552
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 17862 28472 17868 28484
rect 17823 28444 17868 28472
rect 17862 28432 17868 28444
rect 17920 28432 17926 28484
rect 17957 28475 18015 28481
rect 17957 28441 17969 28475
rect 18003 28472 18015 28475
rect 18782 28472 18788 28484
rect 18003 28444 18788 28472
rect 18003 28441 18015 28444
rect 17957 28435 18015 28441
rect 17221 28407 17279 28413
rect 17221 28373 17233 28407
rect 17267 28404 17279 28407
rect 17972 28404 18000 28435
rect 18782 28432 18788 28444
rect 18840 28432 18846 28484
rect 19426 28472 19432 28484
rect 19387 28444 19432 28472
rect 19426 28432 19432 28444
rect 19484 28432 19490 28484
rect 19521 28475 19579 28481
rect 19521 28441 19533 28475
rect 19567 28472 19579 28475
rect 19978 28472 19984 28484
rect 19567 28444 19984 28472
rect 19567 28441 19579 28444
rect 19521 28435 19579 28441
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 20708 28475 20766 28481
rect 20708 28441 20720 28475
rect 20754 28472 20766 28475
rect 21082 28472 21088 28484
rect 20754 28444 21088 28472
rect 20754 28441 20766 28444
rect 20708 28435 20766 28441
rect 21082 28432 21088 28444
rect 21140 28432 21146 28484
rect 22480 28472 22508 28503
rect 21192 28444 22508 28472
rect 18230 28404 18236 28416
rect 17267 28376 18000 28404
rect 18191 28376 18236 28404
rect 17267 28373 17279 28376
rect 17221 28367 17279 28373
rect 18230 28364 18236 28376
rect 18288 28364 18294 28416
rect 20622 28364 20628 28416
rect 20680 28404 20686 28416
rect 21192 28404 21220 28444
rect 21818 28404 21824 28416
rect 20680 28376 21220 28404
rect 21779 28376 21824 28404
rect 20680 28364 20686 28376
rect 21818 28364 21824 28376
rect 21876 28364 21882 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 15841 28203 15899 28209
rect 15841 28169 15853 28203
rect 15887 28200 15899 28203
rect 15930 28200 15936 28212
rect 15887 28172 15936 28200
rect 15887 28169 15899 28172
rect 15841 28163 15899 28169
rect 15930 28160 15936 28172
rect 15988 28160 15994 28212
rect 16850 28160 16856 28212
rect 16908 28200 16914 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16908 28172 17049 28200
rect 16908 28160 16914 28172
rect 17037 28169 17049 28172
rect 17083 28169 17095 28203
rect 17037 28163 17095 28169
rect 17681 28203 17739 28209
rect 17681 28169 17693 28203
rect 17727 28200 17739 28203
rect 17862 28200 17868 28212
rect 17727 28172 17868 28200
rect 17727 28169 17739 28172
rect 17681 28163 17739 28169
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 18046 28160 18052 28212
rect 18104 28200 18110 28212
rect 18877 28203 18935 28209
rect 18877 28200 18889 28203
rect 18104 28172 18889 28200
rect 18104 28160 18110 28172
rect 18877 28169 18889 28172
rect 18923 28169 18935 28203
rect 18877 28163 18935 28169
rect 19242 28160 19248 28212
rect 19300 28160 19306 28212
rect 20622 28200 20628 28212
rect 20583 28172 20628 28200
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 21082 28200 21088 28212
rect 21043 28172 21088 28200
rect 21082 28160 21088 28172
rect 21140 28160 21146 28212
rect 18230 28132 18236 28144
rect 15672 28104 18236 28132
rect 15013 28067 15071 28073
rect 15013 28033 15025 28067
rect 15059 28064 15071 28067
rect 15378 28064 15384 28076
rect 15059 28036 15384 28064
rect 15059 28033 15071 28036
rect 15013 28027 15071 28033
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15672 28073 15700 28104
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 19260 28132 19288 28160
rect 19260 28104 20484 28132
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28033 15715 28067
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 15657 28027 15715 28033
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 18049 28067 18107 28073
rect 18049 28064 18061 28067
rect 17880 28036 18061 28064
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 15473 27999 15531 28005
rect 15473 27996 15485 27999
rect 15344 27968 15485 27996
rect 15344 27956 15350 27968
rect 15473 27965 15485 27968
rect 15519 27965 15531 27999
rect 15473 27959 15531 27965
rect 16669 27999 16727 28005
rect 16669 27965 16681 27999
rect 16715 27996 16727 27999
rect 17586 27996 17592 28008
rect 16715 27968 17592 27996
rect 16715 27965 16727 27968
rect 16669 27959 16727 27965
rect 14829 27931 14887 27937
rect 14829 27897 14841 27931
rect 14875 27928 14887 27931
rect 16684 27928 16712 27959
rect 17586 27956 17592 27968
rect 17644 27956 17650 28008
rect 14875 27900 16712 27928
rect 14875 27897 14887 27900
rect 14829 27891 14887 27897
rect 17880 27860 17908 28036
rect 18049 28033 18061 28036
rect 18095 28033 18107 28067
rect 18049 28027 18107 28033
rect 18156 28036 19196 28064
rect 18156 28008 18184 28036
rect 19168 28008 19196 28036
rect 19242 28024 19248 28076
rect 19300 28064 19306 28076
rect 20073 28067 20131 28073
rect 20073 28064 20085 28067
rect 19300 28036 19345 28064
rect 19444 28036 20085 28064
rect 19300 28024 19306 28036
rect 18138 27996 18144 28008
rect 18099 27968 18144 27996
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 18322 27996 18328 28008
rect 18283 27968 18328 27996
rect 18322 27956 18328 27968
rect 18380 27956 18386 28008
rect 19150 27996 19156 28008
rect 19063 27968 19156 27996
rect 19150 27956 19156 27968
rect 19208 27996 19214 28008
rect 19337 27999 19395 28005
rect 19337 27996 19349 27999
rect 19208 27968 19349 27996
rect 19208 27956 19214 27968
rect 19337 27965 19349 27968
rect 19383 27965 19395 27999
rect 19337 27959 19395 27965
rect 17954 27888 17960 27940
rect 18012 27928 18018 27940
rect 19444 27928 19472 28036
rect 20073 28033 20085 28036
rect 20119 28033 20131 28067
rect 20254 28064 20260 28076
rect 20215 28036 20260 28064
rect 20073 28027 20131 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20456 28073 20484 28104
rect 22664 28104 24532 28132
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 20441 28067 20499 28073
rect 20441 28033 20453 28067
rect 20487 28033 20499 28067
rect 21266 28064 21272 28076
rect 21227 28036 21272 28064
rect 20441 28027 20499 28033
rect 19521 27999 19579 28005
rect 19521 27965 19533 27999
rect 19567 27996 19579 27999
rect 20162 27996 20168 28008
rect 19567 27968 20168 27996
rect 19567 27965 19579 27968
rect 19521 27959 19579 27965
rect 20162 27956 20168 27968
rect 20220 27956 20226 28008
rect 20364 27996 20392 28027
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 21358 28024 21364 28076
rect 21416 28064 21422 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21416 28036 21833 28064
rect 21416 28024 21422 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 22002 28064 22008 28076
rect 21963 28036 22008 28064
rect 21821 28027 21879 28033
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22664 28073 22692 28104
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22152 28036 22661 28064
rect 22152 28024 22158 28036
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 22916 28067 22974 28073
rect 22916 28033 22928 28067
rect 22962 28064 22974 28067
rect 24394 28064 24400 28076
rect 22962 28036 24400 28064
rect 22962 28033 22974 28036
rect 22916 28027 22974 28033
rect 24394 28024 24400 28036
rect 24452 28024 24458 28076
rect 20806 27996 20812 28008
rect 20364 27968 20812 27996
rect 20806 27956 20812 27968
rect 20864 27956 20870 28008
rect 24504 28005 24532 28104
rect 24756 28067 24814 28073
rect 24756 28033 24768 28067
rect 24802 28064 24814 28067
rect 25130 28064 25136 28076
rect 24802 28036 25136 28064
rect 24802 28033 24814 28036
rect 24756 28027 24814 28033
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 24489 27999 24547 28005
rect 24489 27965 24501 27999
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 18012 27900 19472 27928
rect 18012 27888 18018 27900
rect 18782 27860 18788 27872
rect 17880 27832 18788 27860
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 21818 27860 21824 27872
rect 21779 27832 21824 27860
rect 21818 27820 21824 27832
rect 21876 27820 21882 27872
rect 24029 27863 24087 27869
rect 24029 27829 24041 27863
rect 24075 27860 24087 27863
rect 24210 27860 24216 27872
rect 24075 27832 24216 27860
rect 24075 27829 24087 27832
rect 24029 27823 24087 27829
rect 24210 27820 24216 27832
rect 24268 27820 24274 27872
rect 24504 27860 24532 27959
rect 24762 27860 24768 27872
rect 24504 27832 24768 27860
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 25869 27863 25927 27869
rect 25869 27829 25881 27863
rect 25915 27860 25927 27863
rect 26050 27860 26056 27872
rect 25915 27832 26056 27860
rect 25915 27829 25927 27832
rect 25869 27823 25927 27829
rect 26050 27820 26056 27832
rect 26108 27820 26114 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 20254 27616 20260 27668
rect 20312 27656 20318 27668
rect 20441 27659 20499 27665
rect 20441 27656 20453 27659
rect 20312 27628 20453 27656
rect 20312 27616 20318 27628
rect 20441 27625 20453 27628
rect 20487 27625 20499 27659
rect 20441 27619 20499 27625
rect 17221 27591 17279 27597
rect 17221 27557 17233 27591
rect 17267 27588 17279 27591
rect 18138 27588 18144 27600
rect 17267 27560 18144 27588
rect 17267 27557 17279 27560
rect 17221 27551 17279 27557
rect 18138 27548 18144 27560
rect 18196 27548 18202 27600
rect 19245 27591 19303 27597
rect 19245 27557 19257 27591
rect 19291 27588 19303 27591
rect 19426 27588 19432 27600
rect 19291 27560 19432 27588
rect 19291 27557 19303 27560
rect 19245 27551 19303 27557
rect 19426 27548 19432 27560
rect 19484 27548 19490 27600
rect 24394 27588 24400 27600
rect 24355 27560 24400 27588
rect 24394 27548 24400 27560
rect 24452 27548 24458 27600
rect 15470 27480 15476 27532
rect 15528 27520 15534 27532
rect 15933 27523 15991 27529
rect 15933 27520 15945 27523
rect 15528 27492 15945 27520
rect 15528 27480 15534 27492
rect 15933 27489 15945 27492
rect 15979 27489 15991 27523
rect 15933 27483 15991 27489
rect 17034 27480 17040 27532
rect 17092 27520 17098 27532
rect 17865 27523 17923 27529
rect 17865 27520 17877 27523
rect 17092 27492 17877 27520
rect 17092 27480 17098 27492
rect 17865 27489 17877 27492
rect 17911 27489 17923 27523
rect 17865 27483 17923 27489
rect 19334 27480 19340 27532
rect 19392 27520 19398 27532
rect 19797 27523 19855 27529
rect 19797 27520 19809 27523
rect 19392 27492 19809 27520
rect 19392 27480 19398 27492
rect 19797 27489 19809 27492
rect 19843 27489 19855 27523
rect 19797 27483 19855 27489
rect 21085 27523 21143 27529
rect 21085 27489 21097 27523
rect 21131 27520 21143 27523
rect 21818 27520 21824 27532
rect 21131 27492 21824 27520
rect 21131 27489 21143 27492
rect 21085 27483 21143 27489
rect 21818 27480 21824 27492
rect 21876 27480 21882 27532
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 22152 27492 22197 27520
rect 22152 27480 22158 27492
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27452 14151 27455
rect 15746 27452 15752 27464
rect 14139 27424 15752 27452
rect 14139 27421 14151 27424
rect 14093 27415 14151 27421
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 17405 27455 17463 27461
rect 17405 27421 17417 27455
rect 17451 27452 17463 27455
rect 17494 27452 17500 27464
rect 17451 27424 17500 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 13354 27344 13360 27396
rect 13412 27384 13418 27396
rect 14338 27387 14396 27393
rect 14338 27384 14350 27387
rect 13412 27356 14350 27384
rect 13412 27344 13418 27356
rect 14338 27353 14350 27356
rect 14384 27353 14396 27387
rect 15286 27384 15292 27396
rect 14338 27347 14396 27353
rect 14844 27356 15292 27384
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 14844 27316 14872 27356
rect 15286 27344 15292 27356
rect 15344 27384 15350 27396
rect 16224 27384 16252 27415
rect 17494 27412 17500 27424
rect 17552 27412 17558 27464
rect 18046 27412 18052 27464
rect 18104 27452 18110 27464
rect 18141 27455 18199 27461
rect 18141 27452 18153 27455
rect 18104 27424 18153 27452
rect 18104 27412 18110 27424
rect 18141 27421 18153 27424
rect 18187 27421 18199 27455
rect 18141 27415 18199 27421
rect 19150 27412 19156 27464
rect 19208 27452 19214 27464
rect 19705 27455 19763 27461
rect 19705 27452 19717 27455
rect 19208 27424 19717 27452
rect 19208 27412 19214 27424
rect 19705 27421 19717 27424
rect 19751 27452 19763 27455
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 19751 27424 20913 27452
rect 19751 27421 19763 27424
rect 19705 27415 19763 27421
rect 20901 27421 20913 27424
rect 20947 27421 20959 27455
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 20901 27415 20959 27421
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 25222 27452 25228 27464
rect 25183 27424 25228 27452
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 22370 27393 22376 27396
rect 15344 27356 16252 27384
rect 15344 27344 15350 27356
rect 22364 27347 22376 27393
rect 22428 27384 22434 27396
rect 22428 27356 22464 27384
rect 22370 27344 22376 27347
rect 22428 27344 22434 27356
rect 12492 27288 14872 27316
rect 12492 27276 12498 27288
rect 14918 27276 14924 27328
rect 14976 27316 14982 27328
rect 15473 27319 15531 27325
rect 15473 27316 15485 27319
rect 14976 27288 15485 27316
rect 14976 27276 14982 27288
rect 15473 27285 15485 27288
rect 15519 27285 15531 27319
rect 15473 27279 15531 27285
rect 19613 27319 19671 27325
rect 19613 27285 19625 27319
rect 19659 27316 19671 27319
rect 19978 27316 19984 27328
rect 19659 27288 19984 27316
rect 19659 27285 19671 27288
rect 19613 27279 19671 27285
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 20806 27316 20812 27328
rect 20719 27288 20812 27316
rect 20806 27276 20812 27288
rect 20864 27316 20870 27328
rect 21266 27316 21272 27328
rect 20864 27288 21272 27316
rect 20864 27276 20870 27288
rect 21266 27276 21272 27288
rect 21324 27276 21330 27328
rect 22554 27276 22560 27328
rect 22612 27316 22618 27328
rect 23477 27319 23535 27325
rect 23477 27316 23489 27319
rect 22612 27288 23489 27316
rect 22612 27276 22618 27288
rect 23477 27285 23489 27288
rect 23523 27285 23535 27319
rect 25314 27316 25320 27328
rect 25275 27288 25320 27316
rect 23477 27279 23535 27285
rect 25314 27276 25320 27288
rect 25372 27276 25378 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 13354 27112 13360 27124
rect 13315 27084 13360 27112
rect 13354 27072 13360 27084
rect 13412 27072 13418 27124
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17221 27115 17279 27121
rect 17221 27112 17233 27115
rect 16908 27084 17233 27112
rect 16908 27072 16914 27084
rect 17221 27081 17233 27084
rect 17267 27081 17279 27115
rect 17221 27075 17279 27081
rect 19058 27072 19064 27124
rect 19116 27112 19122 27124
rect 19245 27115 19303 27121
rect 19245 27112 19257 27115
rect 19116 27084 19257 27112
rect 19116 27072 19122 27084
rect 19245 27081 19257 27084
rect 19291 27081 19303 27115
rect 19245 27075 19303 27081
rect 20162 27072 20168 27124
rect 20220 27112 20226 27124
rect 20533 27115 20591 27121
rect 20533 27112 20545 27115
rect 20220 27084 20545 27112
rect 20220 27072 20226 27084
rect 20533 27081 20545 27084
rect 20579 27081 20591 27115
rect 20533 27075 20591 27081
rect 15746 27044 15752 27056
rect 14660 27016 15752 27044
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26945 13599 26979
rect 14182 26976 14188 26988
rect 14143 26948 14188 26976
rect 13541 26939 13599 26945
rect 13556 26772 13584 26939
rect 14182 26936 14188 26948
rect 14240 26936 14246 26988
rect 14660 26985 14688 27016
rect 15746 27004 15752 27016
rect 15804 27004 15810 27056
rect 16945 27047 17003 27053
rect 16945 27013 16957 27047
rect 16991 27044 17003 27047
rect 17402 27044 17408 27056
rect 16991 27016 17408 27044
rect 16991 27013 17003 27016
rect 16945 27007 17003 27013
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 17954 27004 17960 27056
rect 18012 27044 18018 27056
rect 18012 27016 18276 27044
rect 18012 27004 18018 27016
rect 14645 26979 14703 26985
rect 14645 26945 14657 26979
rect 14691 26945 14703 26979
rect 14901 26979 14959 26985
rect 14901 26976 14913 26979
rect 14645 26939 14703 26945
rect 14752 26948 14913 26976
rect 14752 26908 14780 26948
rect 14901 26945 14913 26948
rect 14947 26945 14959 26979
rect 14901 26939 14959 26945
rect 16206 26936 16212 26988
rect 16264 26976 16270 26988
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 16264 26948 16681 26976
rect 16264 26936 16270 26948
rect 16669 26945 16681 26948
rect 16715 26945 16727 26979
rect 16850 26976 16856 26988
rect 16811 26948 16856 26976
rect 16669 26939 16727 26945
rect 14016 26880 14780 26908
rect 14016 26849 14044 26880
rect 14001 26843 14059 26849
rect 14001 26809 14013 26843
rect 14047 26809 14059 26843
rect 16684 26840 16712 26939
rect 16850 26936 16856 26948
rect 16908 26936 16914 26988
rect 17034 26976 17040 26988
rect 16995 26948 17040 26976
rect 17034 26936 17040 26948
rect 17092 26936 17098 26988
rect 18248 26985 18276 27016
rect 19150 27004 19156 27056
rect 19208 27044 19214 27056
rect 19705 27047 19763 27053
rect 19705 27044 19717 27047
rect 19208 27016 19717 27044
rect 19208 27004 19214 27016
rect 19705 27013 19717 27016
rect 19751 27013 19763 27047
rect 19705 27007 19763 27013
rect 19794 27004 19800 27056
rect 19852 27044 19858 27056
rect 25222 27044 25228 27056
rect 19852 27016 21312 27044
rect 19852 27004 19858 27016
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 19613 26979 19671 26985
rect 19613 26945 19625 26979
rect 19659 26976 19671 26979
rect 19659 26948 19840 26976
rect 19659 26945 19671 26948
rect 19613 26939 19671 26945
rect 17957 26911 18015 26917
rect 17957 26877 17969 26911
rect 18003 26877 18015 26911
rect 17957 26871 18015 26877
rect 17972 26840 18000 26871
rect 16684 26812 18000 26840
rect 19812 26840 19840 26948
rect 20254 26936 20260 26988
rect 20312 26976 20318 26988
rect 20640 26985 20668 27016
rect 20441 26979 20499 26985
rect 20441 26976 20453 26979
rect 20312 26948 20453 26976
rect 20312 26936 20318 26948
rect 20441 26945 20453 26948
rect 20487 26945 20499 26979
rect 20441 26939 20499 26945
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 20625 26939 20683 26945
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 21284 26985 21312 27016
rect 22112 27016 25228 27044
rect 22112 26985 22140 27016
rect 25222 27004 25228 27016
rect 25280 27044 25286 27056
rect 25501 27047 25559 27053
rect 25280 27016 25360 27044
rect 25280 27004 25286 27016
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20772 26948 21097 26976
rect 20772 26936 20778 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22554 26976 22560 26988
rect 22515 26948 22560 26976
rect 22097 26939 22155 26945
rect 19889 26911 19947 26917
rect 19889 26877 19901 26911
rect 19935 26908 19947 26911
rect 21177 26911 21235 26917
rect 21177 26908 21189 26911
rect 19935 26880 21189 26908
rect 19935 26877 19947 26880
rect 19889 26871 19947 26877
rect 21177 26877 21189 26880
rect 21223 26877 21235 26911
rect 21177 26871 21235 26877
rect 21634 26868 21640 26920
rect 21692 26908 21698 26920
rect 22112 26908 22140 26939
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 25332 26985 25360 27016
rect 25501 27013 25513 27047
rect 25547 27044 25559 27047
rect 26234 27044 26240 27056
rect 25547 27016 26240 27044
rect 25547 27013 25559 27016
rect 25501 27007 25559 27013
rect 26234 27004 26240 27016
rect 26292 27004 26298 27056
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23768 26948 23949 26976
rect 21692 26880 22140 26908
rect 22833 26911 22891 26917
rect 21692 26868 21698 26880
rect 22833 26877 22845 26911
rect 22879 26877 22891 26911
rect 22833 26871 22891 26877
rect 20346 26840 20352 26852
rect 19812 26812 20352 26840
rect 14001 26803 14059 26809
rect 20346 26800 20352 26812
rect 20404 26800 20410 26852
rect 21818 26800 21824 26852
rect 21876 26840 21882 26852
rect 22848 26840 22876 26871
rect 21876 26812 22876 26840
rect 23768 26840 23796 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 24397 26979 24455 26985
rect 24397 26945 24409 26979
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 25317 26979 25375 26985
rect 25317 26945 25329 26979
rect 25363 26945 25375 26979
rect 25317 26939 25375 26945
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26945 25651 26979
rect 26050 26976 26056 26988
rect 26011 26948 26056 26976
rect 25593 26939 25651 26945
rect 23842 26868 23848 26920
rect 23900 26908 23906 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 23900 26880 24133 26908
rect 23900 26868 23906 26880
rect 24121 26877 24133 26880
rect 24167 26877 24179 26911
rect 24121 26871 24179 26877
rect 24210 26868 24216 26920
rect 24268 26908 24274 26920
rect 24412 26908 24440 26939
rect 24762 26908 24768 26920
rect 24268 26880 24313 26908
rect 24412 26880 24768 26908
rect 24268 26868 24274 26880
rect 24762 26868 24768 26880
rect 24820 26908 24826 26920
rect 25608 26908 25636 26939
rect 26050 26936 26056 26948
rect 26108 26936 26114 26988
rect 26878 26936 26884 26988
rect 26936 26976 26942 26988
rect 27229 26979 27287 26985
rect 27229 26976 27241 26979
rect 26936 26948 27241 26976
rect 26936 26936 26942 26948
rect 27229 26945 27241 26948
rect 27275 26945 27287 26979
rect 27229 26939 27287 26945
rect 24820 26880 25636 26908
rect 26973 26911 27031 26917
rect 24820 26868 24826 26880
rect 26973 26877 26985 26911
rect 27019 26877 27031 26911
rect 26973 26871 27031 26877
rect 24026 26840 24032 26852
rect 23768 26812 23888 26840
rect 23987 26812 24032 26840
rect 21876 26800 21882 26812
rect 15930 26772 15936 26784
rect 13556 26744 15936 26772
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 16022 26732 16028 26784
rect 16080 26772 16086 26784
rect 23750 26772 23756 26784
rect 16080 26744 16125 26772
rect 23711 26744 23756 26772
rect 16080 26732 16086 26744
rect 23750 26732 23756 26744
rect 23808 26732 23814 26784
rect 23860 26772 23888 26812
rect 24026 26800 24032 26812
rect 24084 26800 24090 26852
rect 25222 26800 25228 26852
rect 25280 26840 25286 26852
rect 26237 26843 26295 26849
rect 26237 26840 26249 26843
rect 25280 26812 26249 26840
rect 25280 26800 25286 26812
rect 26237 26809 26249 26812
rect 26283 26840 26295 26843
rect 26418 26840 26424 26852
rect 26283 26812 26424 26840
rect 26283 26809 26295 26812
rect 26237 26803 26295 26809
rect 26418 26800 26424 26812
rect 26476 26800 26482 26852
rect 25038 26772 25044 26784
rect 23860 26744 25044 26772
rect 25038 26732 25044 26744
rect 25096 26732 25102 26784
rect 25133 26775 25191 26781
rect 25133 26741 25145 26775
rect 25179 26772 25191 26775
rect 25590 26772 25596 26784
rect 25179 26744 25596 26772
rect 25179 26741 25191 26744
rect 25133 26735 25191 26741
rect 25590 26732 25596 26744
rect 25648 26732 25654 26784
rect 26988 26772 27016 26871
rect 27614 26772 27620 26784
rect 26988 26744 27620 26772
rect 27614 26732 27620 26744
rect 27672 26732 27678 26784
rect 27890 26732 27896 26784
rect 27948 26772 27954 26784
rect 28353 26775 28411 26781
rect 28353 26772 28365 26775
rect 27948 26744 28365 26772
rect 27948 26732 27954 26744
rect 28353 26741 28365 26744
rect 28399 26741 28411 26775
rect 28353 26735 28411 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 14182 26528 14188 26580
rect 14240 26568 14246 26580
rect 15657 26571 15715 26577
rect 15657 26568 15669 26571
rect 14240 26540 15669 26568
rect 14240 26528 14246 26540
rect 15657 26537 15669 26540
rect 15703 26537 15715 26571
rect 15657 26531 15715 26537
rect 15930 26528 15936 26580
rect 15988 26568 15994 26580
rect 16485 26571 16543 26577
rect 16485 26568 16497 26571
rect 15988 26540 16497 26568
rect 15988 26528 15994 26540
rect 16485 26537 16497 26540
rect 16531 26537 16543 26571
rect 16485 26531 16543 26537
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 17037 26571 17095 26577
rect 17037 26568 17049 26571
rect 16908 26540 17049 26568
rect 16908 26528 16914 26540
rect 17037 26537 17049 26540
rect 17083 26537 17095 26571
rect 17037 26531 17095 26537
rect 18322 26528 18328 26580
rect 18380 26568 18386 26580
rect 18509 26571 18567 26577
rect 18509 26568 18521 26571
rect 18380 26540 18521 26568
rect 18380 26528 18386 26540
rect 18509 26537 18521 26540
rect 18555 26537 18567 26571
rect 19334 26568 19340 26580
rect 19295 26540 19340 26568
rect 18509 26531 18567 26537
rect 19334 26528 19340 26540
rect 19392 26528 19398 26580
rect 20898 26528 20904 26580
rect 20956 26568 20962 26580
rect 21269 26571 21327 26577
rect 21269 26568 21281 26571
rect 20956 26540 21281 26568
rect 20956 26528 20962 26540
rect 21269 26537 21281 26540
rect 21315 26537 21327 26571
rect 22186 26568 22192 26580
rect 22147 26540 22192 26568
rect 21269 26531 21327 26537
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 23661 26571 23719 26577
rect 23661 26537 23673 26571
rect 23707 26537 23719 26571
rect 23842 26568 23848 26580
rect 23803 26540 23848 26568
rect 23661 26531 23719 26537
rect 14829 26503 14887 26509
rect 14829 26469 14841 26503
rect 14875 26469 14887 26503
rect 14829 26463 14887 26469
rect 14844 26432 14872 26463
rect 19242 26460 19248 26512
rect 19300 26500 19306 26512
rect 22646 26500 22652 26512
rect 19300 26472 20024 26500
rect 19300 26460 19306 26472
rect 17681 26435 17739 26441
rect 14844 26404 16344 26432
rect 12434 26324 12440 26376
rect 12492 26364 12498 26376
rect 12805 26367 12863 26373
rect 12805 26364 12817 26367
rect 12492 26336 12817 26364
rect 12492 26324 12498 26336
rect 12805 26333 12817 26336
rect 12851 26333 12863 26367
rect 12805 26327 12863 26333
rect 12989 26367 13047 26373
rect 12989 26333 13001 26367
rect 13035 26364 13047 26367
rect 13630 26364 13636 26376
rect 13035 26336 13636 26364
rect 13035 26333 13047 26336
rect 12989 26327 13047 26333
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 14645 26367 14703 26373
rect 14645 26333 14657 26367
rect 14691 26364 14703 26367
rect 15010 26364 15016 26376
rect 14691 26336 15016 26364
rect 14691 26333 14703 26336
rect 14645 26327 14703 26333
rect 13078 26256 13084 26308
rect 13136 26296 13142 26308
rect 14292 26296 14320 26327
rect 15010 26324 15016 26336
rect 15068 26324 15074 26376
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26333 15439 26367
rect 15381 26327 15439 26333
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26364 15531 26367
rect 15930 26364 15936 26376
rect 15519 26336 15936 26364
rect 15519 26333 15531 26336
rect 15473 26327 15531 26333
rect 14458 26296 14464 26308
rect 13136 26268 14320 26296
rect 14419 26268 14464 26296
rect 13136 26256 13142 26268
rect 14458 26256 14464 26268
rect 14516 26256 14522 26308
rect 14553 26299 14611 26305
rect 14553 26265 14565 26299
rect 14599 26296 14611 26299
rect 14918 26296 14924 26308
rect 14599 26268 14924 26296
rect 14599 26265 14611 26268
rect 14553 26259 14611 26265
rect 14918 26256 14924 26268
rect 14976 26256 14982 26308
rect 15396 26296 15424 26327
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16316 26373 16344 26404
rect 17681 26401 17693 26435
rect 17727 26432 17739 26435
rect 19058 26432 19064 26444
rect 17727 26404 19064 26432
rect 17727 26401 17739 26404
rect 17681 26395 17739 26401
rect 19058 26392 19064 26404
rect 19116 26392 19122 26444
rect 16117 26367 16175 26373
rect 16117 26333 16129 26367
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 15654 26296 15660 26308
rect 15396 26268 15660 26296
rect 15654 26256 15660 26268
rect 15712 26296 15718 26308
rect 16132 26296 16160 26327
rect 18230 26324 18236 26376
rect 18288 26364 18294 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18288 26336 18521 26364
rect 18288 26324 18294 26336
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26333 18751 26367
rect 19334 26364 19340 26376
rect 19295 26336 19340 26364
rect 18693 26327 18751 26333
rect 17402 26296 17408 26308
rect 15712 26268 16160 26296
rect 17363 26268 17408 26296
rect 15712 26256 15718 26268
rect 17402 26256 17408 26268
rect 17460 26256 17466 26308
rect 17494 26256 17500 26308
rect 17552 26296 17558 26308
rect 17552 26268 17645 26296
rect 17552 26256 17558 26268
rect 18598 26256 18604 26308
rect 18656 26296 18662 26308
rect 18708 26296 18736 26327
rect 19334 26324 19340 26336
rect 19392 26324 19398 26376
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26364 19579 26367
rect 19794 26364 19800 26376
rect 19567 26336 19800 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 19536 26296 19564 26327
rect 19794 26324 19800 26336
rect 19852 26324 19858 26376
rect 18656 26268 19564 26296
rect 19996 26296 20024 26472
rect 21008 26472 22652 26500
rect 21008 26441 21036 26472
rect 22646 26460 22652 26472
rect 22704 26460 22710 26512
rect 23676 26500 23704 26531
rect 23842 26528 23848 26540
rect 23900 26528 23906 26580
rect 24026 26528 24032 26580
rect 24084 26568 24090 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 24084 26540 24409 26568
rect 24084 26528 24090 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 25130 26568 25136 26580
rect 25091 26540 25136 26568
rect 24397 26531 24455 26537
rect 25130 26528 25136 26540
rect 25188 26528 25194 26580
rect 26878 26568 26884 26580
rect 26839 26540 26884 26568
rect 26878 26528 26884 26540
rect 26936 26528 26942 26580
rect 24210 26500 24216 26512
rect 23676 26472 24216 26500
rect 24210 26460 24216 26472
rect 24268 26500 24274 26512
rect 24268 26472 24716 26500
rect 24268 26460 24274 26472
rect 20993 26435 21051 26441
rect 20993 26401 21005 26435
rect 21039 26401 21051 26435
rect 20993 26395 21051 26401
rect 22005 26435 22063 26441
rect 22005 26401 22017 26435
rect 22051 26432 22063 26435
rect 22051 26404 22600 26432
rect 22051 26401 22063 26404
rect 22005 26395 22063 26401
rect 22572 26376 22600 26404
rect 24688 26376 24716 26472
rect 25222 26460 25228 26512
rect 25280 26500 25286 26512
rect 25501 26503 25559 26509
rect 25501 26500 25513 26503
rect 25280 26472 25513 26500
rect 25280 26460 25286 26472
rect 25501 26469 25513 26472
rect 25547 26500 25559 26503
rect 25547 26472 28212 26500
rect 25547 26469 25559 26472
rect 25501 26463 25559 26469
rect 28184 26441 28212 26472
rect 25409 26435 25467 26441
rect 25409 26401 25421 26435
rect 25455 26432 25467 26435
rect 28169 26435 28227 26441
rect 25455 26404 27108 26432
rect 25455 26401 25467 26404
rect 25409 26395 25467 26401
rect 27080 26376 27108 26404
rect 27172 26404 27927 26432
rect 20073 26367 20131 26373
rect 20073 26333 20085 26367
rect 20119 26364 20131 26367
rect 20162 26364 20168 26376
rect 20119 26336 20168 26364
rect 20119 26333 20131 26336
rect 20073 26327 20131 26333
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20438 26364 20444 26376
rect 20303 26336 20444 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 20901 26367 20959 26373
rect 20901 26333 20913 26367
rect 20947 26364 20959 26367
rect 21634 26364 21640 26376
rect 20947 26336 21640 26364
rect 20947 26333 20959 26336
rect 20901 26327 20959 26333
rect 21634 26324 21640 26336
rect 21692 26324 21698 26376
rect 21913 26367 21971 26373
rect 21913 26333 21925 26367
rect 21959 26364 21971 26367
rect 21959 26336 22094 26364
rect 21959 26333 21971 26336
rect 21913 26327 21971 26333
rect 22066 26296 22094 26336
rect 22554 26324 22560 26376
rect 22612 26364 22618 26376
rect 22741 26367 22799 26373
rect 22741 26364 22753 26367
rect 22612 26336 22753 26364
rect 22612 26324 22618 26336
rect 22741 26333 22753 26336
rect 22787 26333 22799 26367
rect 24670 26364 24676 26376
rect 24631 26336 24676 26364
rect 22741 26327 22799 26333
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 25314 26364 25320 26376
rect 25275 26336 25320 26364
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 25648 26336 25693 26364
rect 25648 26324 25654 26336
rect 25774 26324 25780 26376
rect 25832 26364 25838 26376
rect 26234 26364 26240 26376
rect 25832 26336 25877 26364
rect 26195 26336 26240 26364
rect 25832 26324 25838 26336
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26418 26364 26424 26376
rect 26379 26336 26424 26364
rect 26418 26324 26424 26336
rect 26476 26324 26482 26376
rect 27062 26364 27068 26376
rect 26975 26336 27068 26364
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 27172 26373 27200 26404
rect 27899 26376 27927 26404
rect 28169 26401 28181 26435
rect 28215 26401 28227 26435
rect 28169 26395 28227 26401
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 27341 26367 27399 26373
rect 27341 26333 27353 26367
rect 27387 26333 27399 26367
rect 27341 26327 27399 26333
rect 27433 26367 27491 26373
rect 27433 26333 27445 26367
rect 27479 26364 27491 26367
rect 27706 26364 27712 26376
rect 27479 26336 27712 26364
rect 27479 26333 27491 26336
rect 27433 26327 27491 26333
rect 23106 26296 23112 26308
rect 19996 26268 20300 26296
rect 22066 26268 23112 26296
rect 18656 26256 18662 26268
rect 13170 26228 13176 26240
rect 13131 26200 13176 26228
rect 13170 26188 13176 26200
rect 13228 26188 13234 26240
rect 15286 26188 15292 26240
rect 15344 26228 15350 26240
rect 17512 26228 17540 26256
rect 20272 26237 20300 26268
rect 23106 26256 23112 26268
rect 23164 26256 23170 26308
rect 23477 26299 23535 26305
rect 23477 26265 23489 26299
rect 23523 26296 23535 26299
rect 23566 26296 23572 26308
rect 23523 26268 23572 26296
rect 23523 26265 23535 26268
rect 23477 26259 23535 26265
rect 23566 26256 23572 26268
rect 23624 26256 23630 26308
rect 23693 26299 23751 26305
rect 23693 26265 23705 26299
rect 23739 26296 23751 26299
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 23739 26268 24409 26296
rect 23739 26265 23751 26268
rect 23693 26259 23751 26265
rect 24397 26265 24409 26268
rect 24443 26296 24455 26299
rect 26329 26299 26387 26305
rect 26329 26296 26341 26299
rect 24443 26268 26341 26296
rect 24443 26265 24455 26268
rect 24397 26259 24455 26265
rect 26329 26265 26341 26268
rect 26375 26265 26387 26299
rect 26329 26259 26387 26265
rect 26510 26256 26516 26308
rect 26568 26296 26574 26308
rect 27172 26296 27200 26327
rect 26568 26268 27200 26296
rect 27356 26296 27384 26327
rect 27706 26324 27712 26336
rect 27764 26324 27770 26376
rect 27890 26364 27896 26376
rect 27852 26336 27896 26364
rect 27890 26324 27896 26336
rect 27948 26324 27954 26376
rect 27982 26324 27988 26376
rect 28040 26364 28046 26376
rect 28040 26336 28085 26364
rect 28040 26324 28046 26336
rect 27798 26296 27804 26308
rect 27356 26268 27804 26296
rect 26568 26256 26574 26268
rect 27798 26256 27804 26268
rect 27856 26256 27862 26308
rect 15344 26200 17540 26228
rect 20257 26231 20315 26237
rect 15344 26188 15350 26200
rect 20257 26197 20269 26231
rect 20303 26228 20315 26231
rect 22002 26228 22008 26240
rect 20303 26200 22008 26228
rect 20303 26197 20315 26200
rect 20257 26191 20315 26197
rect 22002 26188 22008 26200
rect 22060 26188 22066 26240
rect 22646 26188 22652 26240
rect 22704 26228 22710 26240
rect 22925 26231 22983 26237
rect 22925 26228 22937 26231
rect 22704 26200 22937 26228
rect 22704 26188 22710 26200
rect 22925 26197 22937 26200
rect 22971 26197 22983 26231
rect 23584 26228 23612 26256
rect 24581 26231 24639 26237
rect 24581 26228 24593 26231
rect 23584 26200 24593 26228
rect 22925 26191 22983 26197
rect 24581 26197 24593 26200
rect 24627 26197 24639 26231
rect 24581 26191 24639 26197
rect 28074 26188 28080 26240
rect 28132 26228 28138 26240
rect 28169 26231 28227 26237
rect 28169 26228 28181 26231
rect 28132 26200 28181 26228
rect 28132 26188 28138 26200
rect 28169 26197 28181 26200
rect 28215 26197 28227 26231
rect 28169 26191 28227 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 14093 26027 14151 26033
rect 14093 25993 14105 26027
rect 14139 26024 14151 26027
rect 14458 26024 14464 26036
rect 14139 25996 14464 26024
rect 14139 25993 14151 25996
rect 14093 25987 14151 25993
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 20070 26024 20076 26036
rect 19444 25996 20076 26024
rect 14553 25959 14611 25965
rect 14553 25925 14565 25959
rect 14599 25956 14611 25959
rect 14734 25956 14740 25968
rect 14599 25928 14740 25956
rect 14599 25925 14611 25928
rect 14553 25919 14611 25925
rect 14734 25916 14740 25928
rect 14792 25916 14798 25968
rect 15930 25916 15936 25968
rect 15988 25956 15994 25968
rect 18690 25956 18696 25968
rect 15988 25928 18696 25956
rect 15988 25916 15994 25928
rect 18690 25916 18696 25928
rect 18748 25916 18754 25968
rect 12250 25848 12256 25900
rect 12308 25888 12314 25900
rect 12417 25891 12475 25897
rect 12417 25888 12429 25891
rect 12308 25860 12429 25888
rect 12308 25848 12314 25860
rect 12417 25857 12429 25860
rect 12463 25857 12475 25891
rect 12417 25851 12475 25857
rect 14461 25891 14519 25897
rect 14461 25857 14473 25891
rect 14507 25888 14519 25891
rect 14918 25888 14924 25900
rect 14507 25860 14924 25888
rect 14507 25857 14519 25860
rect 14461 25851 14519 25857
rect 14918 25848 14924 25860
rect 14976 25848 14982 25900
rect 16850 25888 16856 25900
rect 16811 25860 16856 25888
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25888 17095 25891
rect 17681 25891 17739 25897
rect 17681 25888 17693 25891
rect 17083 25860 17693 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 17681 25857 17693 25860
rect 17727 25857 17739 25891
rect 17681 25851 17739 25857
rect 18417 25891 18475 25897
rect 18417 25857 18429 25891
rect 18463 25857 18475 25891
rect 18598 25888 18604 25900
rect 18559 25860 18604 25888
rect 18417 25851 18475 25857
rect 11790 25780 11796 25832
rect 11848 25820 11854 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 11848 25792 12173 25820
rect 11848 25780 11854 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25789 14795 25823
rect 14737 25783 14795 25789
rect 15289 25823 15347 25829
rect 15289 25789 15301 25823
rect 15335 25820 15347 25823
rect 15470 25820 15476 25832
rect 15335 25792 15476 25820
rect 15335 25789 15347 25792
rect 15289 25783 15347 25789
rect 14752 25752 14780 25783
rect 15470 25780 15476 25792
rect 15528 25780 15534 25832
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25820 15623 25823
rect 15654 25820 15660 25832
rect 15611 25792 15660 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 15654 25780 15660 25792
rect 15712 25820 15718 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 15712 25792 16681 25820
rect 15712 25780 15718 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 18432 25820 18460 25851
rect 18598 25848 18604 25860
rect 18656 25848 18662 25900
rect 19444 25897 19472 25996
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 20993 26027 21051 26033
rect 20993 25993 21005 26027
rect 21039 26024 21051 26027
rect 21358 26024 21364 26036
rect 21039 25996 21364 26024
rect 21039 25993 21051 25996
rect 20993 25987 21051 25993
rect 21008 25956 21036 25987
rect 21358 25984 21364 25996
rect 21416 25984 21422 26036
rect 25314 25984 25320 26036
rect 25372 26024 25378 26036
rect 25372 25996 26464 26024
rect 25372 25984 25378 25996
rect 22738 25956 22744 25968
rect 19812 25928 21036 25956
rect 22020 25928 22744 25956
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25857 19487 25891
rect 19812 25886 19840 25928
rect 19889 25891 19947 25897
rect 19889 25886 19901 25891
rect 19812 25858 19901 25886
rect 19429 25851 19487 25857
rect 19889 25857 19901 25858
rect 19935 25857 19947 25891
rect 20070 25888 20076 25900
rect 20031 25860 20076 25888
rect 19889 25851 19947 25857
rect 18506 25820 18512 25832
rect 18432 25792 18512 25820
rect 16669 25783 16727 25789
rect 18506 25780 18512 25792
rect 18564 25780 18570 25832
rect 19260 25820 19288 25851
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20622 25888 20628 25900
rect 20583 25860 20628 25888
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 20806 25888 20812 25900
rect 20767 25860 20812 25888
rect 20806 25848 20812 25860
rect 20864 25848 20870 25900
rect 22020 25897 22048 25928
rect 22738 25916 22744 25928
rect 22796 25916 22802 25968
rect 26436 25965 26464 25996
rect 27062 25984 27068 26036
rect 27120 26024 27126 26036
rect 27341 26027 27399 26033
rect 27341 26024 27353 26027
rect 27120 25996 27353 26024
rect 27120 25984 27126 25996
rect 27341 25993 27353 25996
rect 27387 26024 27399 26027
rect 27387 25996 27844 26024
rect 27387 25993 27399 25996
rect 27341 25987 27399 25993
rect 27816 25965 27844 25996
rect 24581 25959 24639 25965
rect 24581 25925 24593 25959
rect 24627 25956 24639 25959
rect 26421 25959 26479 25965
rect 24627 25928 25544 25956
rect 24627 25925 24639 25928
rect 24581 25919 24639 25925
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25888 21879 25891
rect 22005 25891 22063 25897
rect 21867 25860 21901 25888
rect 21867 25857 21879 25860
rect 21821 25851 21879 25857
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 20714 25820 20720 25832
rect 19260 25792 20720 25820
rect 20714 25780 20720 25792
rect 20772 25780 20778 25832
rect 21266 25780 21272 25832
rect 21324 25820 21330 25832
rect 21836 25820 21864 25851
rect 22554 25848 22560 25900
rect 22612 25888 22618 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22612 25860 22661 25888
rect 22612 25848 22618 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22830 25888 22836 25900
rect 22791 25860 22836 25888
rect 22649 25851 22707 25857
rect 22830 25848 22836 25860
rect 22888 25848 22894 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 22940 25860 23673 25888
rect 22940 25820 22968 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 24302 25888 24308 25900
rect 24263 25860 24308 25888
rect 23661 25851 23719 25857
rect 24302 25848 24308 25860
rect 24360 25848 24366 25900
rect 24397 25891 24455 25897
rect 24397 25857 24409 25891
rect 24443 25888 24455 25891
rect 25314 25888 25320 25900
rect 24443 25860 25320 25888
rect 24443 25857 24455 25860
rect 24397 25851 24455 25857
rect 21324 25792 22968 25820
rect 21324 25780 21330 25792
rect 23106 25780 23112 25832
rect 23164 25820 23170 25832
rect 24412 25820 24440 25851
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 25516 25897 25544 25928
rect 26421 25925 26433 25959
rect 26467 25956 26479 25959
rect 27801 25959 27859 25965
rect 26467 25928 27292 25956
rect 26467 25925 26479 25928
rect 26421 25919 26479 25925
rect 25409 25891 25467 25897
rect 25409 25857 25421 25891
rect 25455 25857 25467 25891
rect 25409 25851 25467 25857
rect 25501 25891 25559 25897
rect 25501 25857 25513 25891
rect 25547 25857 25559 25891
rect 25501 25851 25559 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25857 25743 25891
rect 26234 25888 26240 25900
rect 26195 25860 26240 25888
rect 25685 25851 25743 25857
rect 23164 25792 24440 25820
rect 24581 25823 24639 25829
rect 23164 25780 23170 25792
rect 24581 25789 24593 25823
rect 24627 25820 24639 25823
rect 24762 25820 24768 25832
rect 24627 25792 24768 25820
rect 24627 25789 24639 25792
rect 24581 25783 24639 25789
rect 24762 25780 24768 25792
rect 24820 25820 24826 25832
rect 25424 25820 25452 25851
rect 24820 25792 25452 25820
rect 24820 25780 24826 25792
rect 19245 25755 19303 25761
rect 19245 25752 19257 25755
rect 14752 25724 19257 25752
rect 19245 25721 19257 25724
rect 19291 25721 19303 25755
rect 19245 25715 19303 25721
rect 25406 25712 25412 25764
rect 25464 25752 25470 25764
rect 25700 25752 25728 25851
rect 26234 25848 26240 25860
rect 26292 25848 26298 25900
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 27264 25888 27292 25928
rect 27801 25925 27813 25959
rect 27847 25925 27859 25959
rect 27801 25919 27859 25925
rect 27985 25959 28043 25965
rect 27985 25925 27997 25959
rect 28031 25956 28043 25959
rect 28626 25956 28632 25968
rect 28031 25928 28632 25956
rect 28031 25925 28043 25928
rect 27985 25919 28043 25925
rect 28626 25916 28632 25928
rect 28684 25916 28690 25968
rect 27890 25888 27896 25900
rect 27264 25860 27896 25888
rect 27890 25848 27896 25860
rect 27948 25848 27954 25900
rect 28074 25848 28080 25900
rect 28132 25888 28138 25900
rect 28132 25860 28177 25888
rect 28132 25848 28138 25860
rect 28258 25848 28264 25900
rect 28316 25888 28322 25900
rect 28537 25891 28595 25897
rect 28537 25888 28549 25891
rect 28316 25860 28549 25888
rect 28316 25848 28322 25860
rect 28537 25857 28549 25860
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25857 28779 25891
rect 28721 25851 28779 25857
rect 26786 25780 26792 25832
rect 26844 25820 26850 25832
rect 26973 25823 27031 25829
rect 26973 25820 26985 25823
rect 26844 25792 26985 25820
rect 26844 25780 26850 25792
rect 26973 25789 26985 25792
rect 27019 25789 27031 25823
rect 26973 25783 27031 25789
rect 27706 25780 27712 25832
rect 27764 25820 27770 25832
rect 28736 25820 28764 25851
rect 30558 25848 30564 25900
rect 30616 25888 30622 25900
rect 31113 25891 31171 25897
rect 31113 25888 31125 25891
rect 30616 25860 31125 25888
rect 30616 25848 30622 25860
rect 31113 25857 31125 25860
rect 31159 25857 31171 25891
rect 31113 25851 31171 25857
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25857 31355 25891
rect 31297 25851 31355 25857
rect 27764 25792 28764 25820
rect 27764 25780 27770 25792
rect 29362 25780 29368 25832
rect 29420 25820 29426 25832
rect 31312 25820 31340 25851
rect 34790 25820 34796 25832
rect 29420 25792 34796 25820
rect 29420 25780 29426 25792
rect 34790 25780 34796 25792
rect 34848 25780 34854 25832
rect 27798 25752 27804 25764
rect 25464 25724 25728 25752
rect 27759 25724 27804 25752
rect 25464 25712 25470 25724
rect 27798 25712 27804 25724
rect 27856 25712 27862 25764
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 13541 25687 13599 25693
rect 13541 25684 13553 25687
rect 13320 25656 13553 25684
rect 13320 25644 13326 25656
rect 13541 25653 13553 25656
rect 13587 25653 13599 25687
rect 17494 25684 17500 25696
rect 17455 25656 17500 25684
rect 13541 25647 13599 25653
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 18414 25684 18420 25696
rect 18375 25656 18420 25684
rect 18414 25644 18420 25656
rect 18472 25644 18478 25696
rect 19886 25684 19892 25696
rect 19847 25656 19892 25684
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 20809 25687 20867 25693
rect 20809 25653 20821 25687
rect 20855 25684 20867 25687
rect 20898 25684 20904 25696
rect 20855 25656 20904 25684
rect 20855 25653 20867 25656
rect 20809 25647 20867 25653
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 21913 25687 21971 25693
rect 21913 25653 21925 25687
rect 21959 25684 21971 25687
rect 22462 25684 22468 25696
rect 21959 25656 22468 25684
rect 21959 25653 21971 25656
rect 21913 25647 21971 25653
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 25041 25687 25099 25693
rect 25041 25653 25053 25687
rect 25087 25684 25099 25687
rect 25682 25684 25688 25696
rect 25087 25656 25688 25684
rect 25087 25653 25099 25656
rect 25041 25647 25099 25653
rect 25682 25644 25688 25656
rect 25740 25644 25746 25696
rect 27890 25644 27896 25696
rect 27948 25684 27954 25696
rect 28537 25687 28595 25693
rect 28537 25684 28549 25687
rect 27948 25656 28549 25684
rect 27948 25644 27954 25656
rect 28537 25653 28549 25656
rect 28583 25653 28595 25687
rect 28537 25647 28595 25653
rect 31205 25687 31263 25693
rect 31205 25653 31217 25687
rect 31251 25684 31263 25687
rect 32858 25684 32864 25696
rect 31251 25656 32864 25684
rect 31251 25653 31263 25656
rect 31205 25647 31263 25653
rect 32858 25644 32864 25656
rect 32916 25644 32922 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 12161 25483 12219 25489
rect 12161 25449 12173 25483
rect 12207 25480 12219 25483
rect 12250 25480 12256 25492
rect 12207 25452 12256 25480
rect 12207 25449 12219 25452
rect 12161 25443 12219 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 19886 25480 19892 25492
rect 13464 25452 19892 25480
rect 5258 25304 5264 25356
rect 5316 25344 5322 25356
rect 13464 25353 13492 25452
rect 19886 25440 19892 25452
rect 19944 25440 19950 25492
rect 20533 25483 20591 25489
rect 20533 25449 20545 25483
rect 20579 25480 20591 25483
rect 20898 25480 20904 25492
rect 20579 25452 20904 25480
rect 20579 25449 20591 25452
rect 20533 25443 20591 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 23845 25483 23903 25489
rect 23845 25449 23857 25483
rect 23891 25480 23903 25483
rect 24578 25480 24584 25492
rect 23891 25452 24584 25480
rect 23891 25449 23903 25452
rect 23845 25443 23903 25449
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 24762 25440 24768 25492
rect 24820 25480 24826 25492
rect 25041 25483 25099 25489
rect 25041 25480 25053 25483
rect 24820 25452 25053 25480
rect 24820 25440 24826 25452
rect 25041 25449 25053 25452
rect 25087 25449 25099 25483
rect 25041 25443 25099 25449
rect 18046 25372 18052 25424
rect 18104 25412 18110 25424
rect 19245 25415 19303 25421
rect 19245 25412 19257 25415
rect 18104 25384 19257 25412
rect 18104 25372 18110 25384
rect 19245 25381 19257 25384
rect 19291 25381 19303 25415
rect 20714 25412 20720 25424
rect 20675 25384 20720 25412
rect 19245 25375 19303 25381
rect 20714 25372 20720 25384
rect 20772 25372 20778 25424
rect 21266 25412 21272 25424
rect 21100 25384 21272 25412
rect 13449 25347 13507 25353
rect 5316 25316 13400 25344
rect 5316 25304 5322 25316
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 13170 25276 13176 25288
rect 12391 25248 13176 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 13170 25236 13176 25248
rect 13228 25236 13234 25288
rect 13372 25276 13400 25316
rect 13449 25313 13461 25347
rect 13495 25313 13507 25347
rect 15286 25344 15292 25356
rect 13449 25307 13507 25313
rect 14660 25316 15292 25344
rect 14660 25285 14688 25316
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 15746 25304 15752 25356
rect 15804 25344 15810 25356
rect 16298 25344 16304 25356
rect 15804 25316 16304 25344
rect 15804 25304 15810 25316
rect 16298 25304 16304 25316
rect 16356 25304 16362 25356
rect 20254 25344 20260 25356
rect 19260 25316 20260 25344
rect 14645 25279 14703 25285
rect 14645 25276 14657 25279
rect 13372 25248 14657 25276
rect 14645 25245 14657 25248
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 14734 25236 14740 25288
rect 14792 25276 14798 25288
rect 14921 25279 14979 25285
rect 14921 25276 14933 25279
rect 14792 25248 14933 25276
rect 14792 25236 14798 25248
rect 14921 25245 14933 25248
rect 14967 25245 14979 25279
rect 14921 25239 14979 25245
rect 16568 25279 16626 25285
rect 16568 25245 16580 25279
rect 16614 25276 16626 25279
rect 17494 25276 17500 25288
rect 16614 25248 17500 25276
rect 16614 25245 16626 25248
rect 16568 25239 16626 25245
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 18230 25276 18236 25288
rect 18191 25248 18236 25276
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 19260 25285 19288 25316
rect 20254 25304 20260 25316
rect 20312 25304 20318 25356
rect 20441 25347 20499 25353
rect 20441 25313 20453 25347
rect 20487 25344 20499 25347
rect 21100 25344 21128 25384
rect 21266 25372 21272 25384
rect 21324 25372 21330 25424
rect 20487 25316 21128 25344
rect 21177 25347 21235 25353
rect 20487 25313 20499 25316
rect 20441 25307 20499 25313
rect 21177 25313 21189 25347
rect 21223 25344 21235 25347
rect 22462 25344 22468 25356
rect 21223 25316 22468 25344
rect 21223 25313 21235 25316
rect 21177 25307 21235 25313
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 22554 25304 22560 25356
rect 22612 25344 22618 25356
rect 23014 25344 23020 25356
rect 22612 25316 22657 25344
rect 22975 25316 23020 25344
rect 22612 25304 22618 25316
rect 23014 25304 23020 25316
rect 23072 25304 23078 25356
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 25593 25347 25651 25353
rect 25593 25344 25605 25347
rect 24912 25316 25605 25344
rect 24912 25304 24918 25316
rect 25593 25313 25605 25316
rect 25639 25313 25651 25347
rect 25593 25307 25651 25313
rect 19426 25285 19432 25288
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 19423 25276 19432 25285
rect 19245 25239 19303 25245
rect 19352 25248 19432 25276
rect 13265 25211 13323 25217
rect 13265 25177 13277 25211
rect 13311 25208 13323 25211
rect 14752 25208 14780 25236
rect 13311 25180 14780 25208
rect 18432 25208 18460 25239
rect 19352 25208 19380 25248
rect 19423 25239 19432 25248
rect 19426 25236 19432 25239
rect 19484 25236 19490 25288
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25245 20407 25279
rect 20349 25239 20407 25245
rect 18432 25180 19380 25208
rect 20364 25208 20392 25239
rect 20806 25236 20812 25288
rect 20864 25276 20870 25288
rect 21453 25279 21511 25285
rect 21453 25276 21465 25279
rect 20864 25248 21465 25276
rect 20864 25236 20870 25248
rect 21453 25245 21465 25248
rect 21499 25245 21511 25279
rect 21453 25239 21511 25245
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25276 22707 25279
rect 23106 25276 23112 25288
rect 22695 25248 23112 25276
rect 22695 25245 22707 25248
rect 22649 25239 22707 25245
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25276 23535 25279
rect 23750 25276 23756 25288
rect 23523 25248 23756 25276
rect 23523 25245 23535 25248
rect 23477 25239 23535 25245
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25245 25007 25279
rect 25130 25276 25136 25288
rect 25091 25248 25136 25276
rect 24949 25239 25007 25245
rect 20714 25208 20720 25220
rect 20364 25180 20720 25208
rect 13311 25177 13323 25180
rect 13265 25171 13323 25177
rect 20714 25168 20720 25180
rect 20772 25168 20778 25220
rect 23661 25211 23719 25217
rect 23661 25177 23673 25211
rect 23707 25208 23719 25211
rect 23934 25208 23940 25220
rect 23707 25180 23940 25208
rect 23707 25177 23719 25180
rect 23661 25171 23719 25177
rect 23934 25168 23940 25180
rect 23992 25168 23998 25220
rect 24964 25208 24992 25239
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25682 25236 25688 25288
rect 25740 25276 25746 25288
rect 25849 25279 25907 25285
rect 25849 25276 25861 25279
rect 25740 25248 25861 25276
rect 25740 25236 25746 25248
rect 25849 25245 25861 25248
rect 25895 25245 25907 25279
rect 27614 25276 27620 25288
rect 27575 25248 27620 25276
rect 25849 25239 25907 25245
rect 27614 25236 27620 25248
rect 27672 25236 27678 25288
rect 27890 25285 27896 25288
rect 27884 25276 27896 25285
rect 27851 25248 27896 25276
rect 27884 25239 27896 25248
rect 27890 25236 27896 25239
rect 27948 25236 27954 25288
rect 29822 25276 29828 25288
rect 29783 25248 29828 25276
rect 29822 25236 29828 25248
rect 29880 25276 29886 25288
rect 31662 25276 31668 25288
rect 29880 25248 31668 25276
rect 29880 25236 29886 25248
rect 31662 25236 31668 25248
rect 31720 25236 31726 25288
rect 25038 25208 25044 25220
rect 24951 25180 25044 25208
rect 25038 25168 25044 25180
rect 25096 25208 25102 25220
rect 27154 25208 27160 25220
rect 25096 25180 27160 25208
rect 25096 25168 25102 25180
rect 27154 25168 27160 25180
rect 27212 25168 27218 25220
rect 30092 25211 30150 25217
rect 30092 25177 30104 25211
rect 30138 25208 30150 25211
rect 30466 25208 30472 25220
rect 30138 25180 30472 25208
rect 30138 25177 30150 25180
rect 30092 25171 30150 25177
rect 30466 25168 30472 25180
rect 30524 25168 30530 25220
rect 30742 25168 30748 25220
rect 30800 25208 30806 25220
rect 31910 25211 31968 25217
rect 31910 25208 31922 25211
rect 30800 25180 31922 25208
rect 30800 25168 30806 25180
rect 31910 25177 31922 25180
rect 31956 25177 31968 25211
rect 31910 25171 31968 25177
rect 12802 25140 12808 25152
rect 12763 25112 12808 25140
rect 12802 25100 12808 25112
rect 12860 25100 12866 25152
rect 13170 25140 13176 25152
rect 13131 25112 13176 25140
rect 13170 25100 13176 25112
rect 13228 25100 13234 25152
rect 17218 25100 17224 25152
rect 17276 25140 17282 25152
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17276 25112 17693 25140
rect 17276 25100 17282 25112
rect 17681 25109 17693 25112
rect 17727 25109 17739 25143
rect 17681 25103 17739 25109
rect 17954 25100 17960 25152
rect 18012 25140 18018 25152
rect 18325 25143 18383 25149
rect 18325 25140 18337 25143
rect 18012 25112 18337 25140
rect 18012 25100 18018 25112
rect 18325 25109 18337 25112
rect 18371 25109 18383 25143
rect 18325 25103 18383 25109
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26973 25143 27031 25149
rect 26973 25140 26985 25143
rect 26292 25112 26985 25140
rect 26292 25100 26298 25112
rect 26973 25109 26985 25112
rect 27019 25109 27031 25143
rect 26973 25103 27031 25109
rect 28166 25100 28172 25152
rect 28224 25140 28230 25152
rect 28997 25143 29055 25149
rect 28997 25140 29009 25143
rect 28224 25112 29009 25140
rect 28224 25100 28230 25112
rect 28997 25109 29009 25112
rect 29043 25109 29055 25143
rect 31202 25140 31208 25152
rect 31163 25112 31208 25140
rect 28997 25103 29055 25109
rect 31202 25100 31208 25112
rect 31260 25100 31266 25152
rect 31294 25100 31300 25152
rect 31352 25140 31358 25152
rect 33045 25143 33103 25149
rect 33045 25140 33057 25143
rect 31352 25112 33057 25140
rect 31352 25100 31358 25112
rect 33045 25109 33057 25112
rect 33091 25109 33103 25143
rect 33045 25103 33103 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 17313 24939 17371 24945
rect 17313 24936 17325 24939
rect 17276 24908 17325 24936
rect 17276 24896 17282 24908
rect 17313 24905 17325 24908
rect 17359 24905 17371 24939
rect 18690 24936 18696 24948
rect 18651 24908 18696 24936
rect 17313 24899 17371 24905
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 22051 24939 22109 24945
rect 22051 24905 22063 24939
rect 22097 24905 22109 24939
rect 22051 24899 22109 24905
rect 12802 24828 12808 24880
rect 12860 24868 12866 24880
rect 13265 24871 13323 24877
rect 13265 24868 13277 24871
rect 12860 24840 13277 24868
rect 12860 24828 12866 24840
rect 13265 24837 13277 24840
rect 13311 24837 13323 24871
rect 13265 24831 13323 24837
rect 14461 24871 14519 24877
rect 14461 24837 14473 24871
rect 14507 24868 14519 24871
rect 15194 24868 15200 24880
rect 14507 24840 15200 24868
rect 14507 24837 14519 24840
rect 14461 24831 14519 24837
rect 15194 24828 15200 24840
rect 15252 24828 15258 24880
rect 17236 24840 17448 24868
rect 13078 24800 13084 24812
rect 13039 24772 13084 24800
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 13449 24803 13507 24809
rect 13449 24769 13461 24803
rect 13495 24769 13507 24803
rect 17236 24800 17264 24840
rect 13449 24763 13507 24769
rect 14752 24772 17264 24800
rect 17420 24800 17448 24840
rect 17862 24828 17868 24880
rect 17920 24868 17926 24880
rect 22066 24868 22094 24899
rect 23750 24896 23756 24948
rect 23808 24936 23814 24948
rect 25130 24936 25136 24948
rect 23808 24908 25136 24936
rect 23808 24896 23814 24908
rect 25130 24896 25136 24908
rect 25188 24936 25194 24948
rect 25188 24908 26004 24936
rect 25188 24896 25194 24908
rect 17920 24840 18184 24868
rect 17920 24828 17926 24840
rect 18046 24800 18052 24812
rect 17420 24772 18052 24800
rect 13262 24692 13268 24744
rect 13320 24732 13326 24744
rect 13372 24732 13400 24763
rect 13320 24704 13400 24732
rect 13320 24692 13326 24704
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 13464 24596 13492 24763
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 14642 24732 14648 24744
rect 14599 24704 14648 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14752 24741 14780 24772
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18156 24809 18184 24840
rect 21744 24840 22094 24868
rect 25148 24840 25360 24868
rect 18141 24803 18199 24809
rect 18141 24769 18153 24803
rect 18187 24769 18199 24803
rect 18141 24763 18199 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24701 14795 24735
rect 15286 24732 15292 24744
rect 15247 24704 15292 24732
rect 14737 24695 14795 24701
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 15565 24735 15623 24741
rect 15565 24701 15577 24735
rect 15611 24732 15623 24735
rect 17126 24732 17132 24744
rect 15611 24704 17132 24732
rect 15611 24701 15623 24704
rect 15565 24695 15623 24701
rect 17126 24692 17132 24704
rect 17184 24732 17190 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 17184 24704 17417 24732
rect 17184 24692 17190 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24732 17647 24735
rect 17954 24732 17960 24744
rect 17635 24704 17960 24732
rect 17635 24701 17647 24704
rect 17589 24695 17647 24701
rect 17954 24692 17960 24704
rect 18012 24692 18018 24744
rect 13630 24664 13636 24676
rect 13591 24636 13636 24664
rect 13630 24624 13636 24636
rect 13688 24624 13694 24676
rect 14093 24667 14151 24673
rect 14093 24633 14105 24667
rect 14139 24664 14151 24667
rect 18340 24664 18368 24763
rect 18432 24732 18460 24763
rect 18506 24760 18512 24812
rect 18564 24800 18570 24812
rect 19613 24803 19671 24809
rect 18564 24772 18609 24800
rect 18564 24760 18570 24772
rect 19613 24769 19625 24803
rect 19659 24800 19671 24803
rect 19978 24800 19984 24812
rect 19659 24772 19984 24800
rect 19659 24769 19671 24772
rect 19613 24763 19671 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20622 24800 20628 24812
rect 20535 24772 20628 24800
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20806 24800 20812 24812
rect 20767 24772 20812 24800
rect 20806 24760 20812 24772
rect 20864 24760 20870 24812
rect 21542 24760 21548 24812
rect 21600 24800 21606 24812
rect 21744 24800 21772 24840
rect 21600 24772 21772 24800
rect 21821 24803 21879 24809
rect 21600 24760 21606 24772
rect 21821 24769 21833 24803
rect 21867 24800 21879 24803
rect 23014 24800 23020 24812
rect 21867 24772 23020 24800
rect 21867 24769 21879 24772
rect 21821 24763 21879 24769
rect 23014 24760 23020 24772
rect 23072 24800 23078 24812
rect 23109 24803 23167 24809
rect 23109 24800 23121 24803
rect 23072 24772 23121 24800
rect 23072 24760 23078 24772
rect 23109 24769 23121 24772
rect 23155 24769 23167 24803
rect 24210 24800 24216 24812
rect 24171 24772 24216 24800
rect 23109 24763 23167 24769
rect 24210 24760 24216 24772
rect 24268 24760 24274 24812
rect 24302 24760 24308 24812
rect 24360 24800 24366 24812
rect 24762 24800 24768 24812
rect 24360 24772 24768 24800
rect 24360 24760 24366 24772
rect 24762 24760 24768 24772
rect 24820 24800 24826 24812
rect 25148 24800 25176 24840
rect 24820 24772 25176 24800
rect 25225 24803 25283 24809
rect 24820 24760 24826 24772
rect 25225 24769 25237 24803
rect 25271 24769 25283 24803
rect 25332 24800 25360 24840
rect 25409 24803 25467 24809
rect 25409 24800 25421 24803
rect 25332 24772 25421 24800
rect 25225 24763 25283 24769
rect 25409 24769 25421 24772
rect 25455 24769 25467 24803
rect 25976 24800 26004 24908
rect 26234 24896 26240 24948
rect 26292 24945 26298 24948
rect 26292 24939 26311 24945
rect 26299 24905 26311 24939
rect 26292 24899 26311 24905
rect 26292 24896 26298 24899
rect 27614 24896 27620 24948
rect 27672 24896 27678 24948
rect 27801 24939 27859 24945
rect 27801 24905 27813 24939
rect 27847 24936 27859 24939
rect 28445 24939 28503 24945
rect 28445 24936 28457 24939
rect 27847 24908 28457 24936
rect 27847 24905 27859 24908
rect 27801 24899 27859 24905
rect 28445 24905 28457 24908
rect 28491 24905 28503 24939
rect 28445 24899 28503 24905
rect 26053 24871 26111 24877
rect 26053 24837 26065 24871
rect 26099 24868 26111 24871
rect 26142 24868 26148 24880
rect 26099 24840 26148 24868
rect 26099 24837 26111 24840
rect 26053 24831 26111 24837
rect 26142 24828 26148 24840
rect 26200 24828 26206 24880
rect 27632 24868 27660 24896
rect 29822 24868 29828 24880
rect 27632 24840 29828 24868
rect 26234 24800 26240 24812
rect 25976 24772 26240 24800
rect 25409 24763 25467 24769
rect 18874 24732 18880 24744
rect 18432 24704 18880 24732
rect 18874 24692 18880 24704
rect 18932 24692 18938 24744
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 19337 24735 19395 24741
rect 19337 24732 19349 24735
rect 19300 24704 19349 24732
rect 19300 24692 19306 24704
rect 19337 24701 19349 24704
rect 19383 24701 19395 24735
rect 20640 24732 20668 24760
rect 21910 24732 21916 24744
rect 20640 24704 21916 24732
rect 19337 24695 19395 24701
rect 21910 24692 21916 24704
rect 21968 24692 21974 24744
rect 22462 24692 22468 24744
rect 22520 24732 22526 24744
rect 23201 24735 23259 24741
rect 23201 24732 23213 24735
rect 22520 24704 23213 24732
rect 22520 24692 22526 24704
rect 23201 24701 23213 24704
rect 23247 24701 23259 24735
rect 25240 24732 25268 24763
rect 26234 24760 26240 24772
rect 26292 24800 26298 24812
rect 26786 24800 26792 24812
rect 26292 24772 26792 24800
rect 26292 24760 26298 24772
rect 26786 24760 26792 24772
rect 26844 24760 26850 24812
rect 26970 24800 26976 24812
rect 26931 24772 26976 24800
rect 26970 24760 26976 24772
rect 27028 24760 27034 24812
rect 27617 24803 27675 24809
rect 27617 24769 27629 24803
rect 27663 24800 27675 24803
rect 27706 24800 27712 24812
rect 27663 24772 27712 24800
rect 27663 24769 27675 24772
rect 27617 24763 27675 24769
rect 25590 24732 25596 24744
rect 25240 24704 25596 24732
rect 23201 24695 23259 24701
rect 25590 24692 25596 24704
rect 25648 24732 25654 24744
rect 25648 24704 26372 24732
rect 25648 24692 25654 24704
rect 26344 24676 26372 24704
rect 14139 24636 18368 24664
rect 18984 24636 20760 24664
rect 14139 24633 14151 24636
rect 14093 24627 14151 24633
rect 15010 24596 15016 24608
rect 13412 24568 15016 24596
rect 13412 24556 13418 24568
rect 15010 24556 15016 24568
rect 15068 24556 15074 24608
rect 16945 24599 17003 24605
rect 16945 24565 16957 24599
rect 16991 24596 17003 24599
rect 17494 24596 17500 24608
rect 16991 24568 17500 24596
rect 16991 24565 17003 24568
rect 16945 24559 17003 24565
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 18230 24556 18236 24608
rect 18288 24596 18294 24608
rect 18984 24596 19012 24636
rect 20622 24596 20628 24608
rect 18288 24568 19012 24596
rect 20583 24568 20628 24596
rect 18288 24556 18294 24568
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 20732 24596 20760 24636
rect 20898 24624 20904 24676
rect 20956 24664 20962 24676
rect 20956 24636 22094 24664
rect 20956 24624 20962 24636
rect 20993 24599 21051 24605
rect 20993 24596 21005 24599
rect 20732 24568 21005 24596
rect 20993 24565 21005 24568
rect 21039 24565 21051 24599
rect 22066 24596 22094 24636
rect 22830 24624 22836 24676
rect 22888 24664 22894 24676
rect 25222 24664 25228 24676
rect 22888 24636 25084 24664
rect 25183 24636 25228 24664
rect 22888 24624 22894 24636
rect 23109 24599 23167 24605
rect 23109 24596 23121 24599
rect 22066 24568 23121 24596
rect 20993 24559 21051 24565
rect 23109 24565 23121 24568
rect 23155 24565 23167 24599
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23109 24559 23167 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 24026 24596 24032 24608
rect 23987 24568 24032 24596
rect 24026 24556 24032 24568
rect 24084 24556 24090 24608
rect 25056 24596 25084 24636
rect 25222 24624 25228 24636
rect 25280 24624 25286 24676
rect 26326 24624 26332 24676
rect 26384 24664 26390 24676
rect 26421 24667 26479 24673
rect 26421 24664 26433 24667
rect 26384 24636 26433 24664
rect 26384 24624 26390 24636
rect 26421 24633 26433 24636
rect 26467 24633 26479 24667
rect 27632 24664 27660 24763
rect 27706 24760 27712 24772
rect 27764 24760 27770 24812
rect 27893 24803 27951 24809
rect 27893 24769 27905 24803
rect 27939 24800 27951 24803
rect 27982 24800 27988 24812
rect 27939 24772 27988 24800
rect 27939 24769 27951 24772
rect 27893 24763 27951 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28353 24803 28411 24809
rect 28353 24800 28365 24803
rect 28276 24772 28365 24800
rect 27890 24664 27896 24676
rect 27632 24636 27896 24664
rect 26421 24627 26479 24633
rect 27890 24624 27896 24636
rect 27948 24624 27954 24676
rect 26237 24599 26295 24605
rect 26237 24596 26249 24599
rect 25056 24568 26249 24596
rect 26237 24565 26249 24568
rect 26283 24596 26295 24599
rect 26510 24596 26516 24608
rect 26283 24568 26516 24596
rect 26283 24565 26295 24568
rect 26237 24559 26295 24565
rect 26510 24556 26516 24568
rect 26568 24556 26574 24608
rect 27062 24596 27068 24608
rect 27023 24568 27068 24596
rect 27062 24556 27068 24568
rect 27120 24556 27126 24608
rect 27617 24599 27675 24605
rect 27617 24565 27629 24599
rect 27663 24596 27675 24599
rect 27706 24596 27712 24608
rect 27663 24568 27712 24596
rect 27663 24565 27675 24568
rect 27617 24559 27675 24565
rect 27706 24556 27712 24568
rect 27764 24556 27770 24608
rect 28276 24596 28304 24772
rect 28353 24769 28365 24772
rect 28399 24769 28411 24803
rect 28353 24763 28411 24769
rect 28534 24760 28540 24812
rect 28592 24800 28598 24812
rect 29104 24809 29132 24840
rect 29822 24828 29828 24840
rect 29880 24828 29886 24880
rect 29089 24803 29147 24809
rect 28592 24772 28637 24800
rect 28592 24760 28598 24772
rect 29089 24769 29101 24803
rect 29135 24769 29147 24803
rect 29089 24763 29147 24769
rect 29356 24803 29414 24809
rect 29356 24769 29368 24803
rect 29402 24800 29414 24803
rect 30374 24800 30380 24812
rect 29402 24772 30380 24800
rect 29402 24769 29414 24772
rect 29356 24763 29414 24769
rect 30374 24760 30380 24772
rect 30432 24760 30438 24812
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24769 31079 24803
rect 31021 24763 31079 24769
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24800 32643 24803
rect 32674 24800 32680 24812
rect 32631 24772 32680 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 31036 24732 31064 24763
rect 32674 24760 32680 24772
rect 32732 24760 32738 24812
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 30208 24704 31064 24732
rect 28994 24596 29000 24608
rect 28276 24568 29000 24596
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29822 24556 29828 24608
rect 29880 24596 29886 24608
rect 30208 24596 30236 24704
rect 32030 24692 32036 24744
rect 32088 24732 32094 24744
rect 32784 24732 32812 24763
rect 32088 24704 32812 24732
rect 32088 24692 32094 24704
rect 30282 24624 30288 24676
rect 30340 24664 30346 24676
rect 31205 24667 31263 24673
rect 31205 24664 31217 24667
rect 30340 24636 31217 24664
rect 30340 24624 30346 24636
rect 31205 24633 31217 24636
rect 31251 24633 31263 24667
rect 31205 24627 31263 24633
rect 30469 24599 30527 24605
rect 30469 24596 30481 24599
rect 29880 24568 30481 24596
rect 29880 24556 29886 24568
rect 30469 24565 30481 24568
rect 30515 24565 30527 24599
rect 30469 24559 30527 24565
rect 32306 24556 32312 24608
rect 32364 24596 32370 24608
rect 32585 24599 32643 24605
rect 32585 24596 32597 24599
rect 32364 24568 32597 24596
rect 32364 24556 32370 24568
rect 32585 24565 32597 24568
rect 32631 24565 32643 24599
rect 32585 24559 32643 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 16850 24352 16856 24404
rect 16908 24392 16914 24404
rect 17865 24395 17923 24401
rect 17865 24392 17877 24395
rect 16908 24364 17877 24392
rect 16908 24352 16914 24364
rect 17865 24361 17877 24364
rect 17911 24361 17923 24395
rect 17865 24355 17923 24361
rect 20622 24352 20628 24404
rect 20680 24392 20686 24404
rect 20717 24395 20775 24401
rect 20717 24392 20729 24395
rect 20680 24364 20729 24392
rect 20680 24352 20686 24364
rect 20717 24361 20729 24364
rect 20763 24392 20775 24395
rect 21818 24392 21824 24404
rect 20763 24364 21824 24392
rect 20763 24361 20775 24364
rect 20717 24355 20775 24361
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 24210 24352 24216 24404
rect 24268 24392 24274 24404
rect 24857 24395 24915 24401
rect 24857 24392 24869 24395
rect 24268 24364 24869 24392
rect 24268 24352 24274 24364
rect 24857 24361 24869 24364
rect 24903 24392 24915 24395
rect 25593 24395 25651 24401
rect 25593 24392 25605 24395
rect 24903 24364 25605 24392
rect 24903 24361 24915 24364
rect 24857 24355 24915 24361
rect 25593 24361 25605 24364
rect 25639 24361 25651 24395
rect 25593 24355 25651 24361
rect 26234 24352 26240 24404
rect 26292 24392 26298 24404
rect 26329 24395 26387 24401
rect 26329 24392 26341 24395
rect 26292 24364 26341 24392
rect 26292 24352 26298 24364
rect 26329 24361 26341 24364
rect 26375 24361 26387 24395
rect 26329 24355 26387 24361
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 30009 24395 30067 24401
rect 27856 24364 28396 24392
rect 27856 24352 27862 24364
rect 15194 24284 15200 24336
rect 15252 24324 15258 24336
rect 16022 24324 16028 24336
rect 15252 24296 16028 24324
rect 15252 24284 15258 24296
rect 16022 24284 16028 24296
rect 16080 24324 16086 24336
rect 16080 24296 17816 24324
rect 16080 24284 16086 24296
rect 15010 24256 15016 24268
rect 14971 24228 15016 24256
rect 15010 24216 15016 24228
rect 15068 24216 15074 24268
rect 17788 24256 17816 24296
rect 18322 24284 18328 24336
rect 18380 24324 18386 24336
rect 19245 24327 19303 24333
rect 19245 24324 19257 24327
rect 18380 24296 19257 24324
rect 18380 24284 18386 24296
rect 19245 24293 19257 24296
rect 19291 24293 19303 24327
rect 20901 24327 20959 24333
rect 20901 24324 20913 24327
rect 19245 24287 19303 24293
rect 19352 24296 20913 24324
rect 19352 24268 19380 24296
rect 20901 24293 20913 24296
rect 20947 24293 20959 24327
rect 28368 24324 28396 24364
rect 30009 24361 30021 24395
rect 30055 24392 30067 24395
rect 30055 24364 30696 24392
rect 30055 24361 30067 24364
rect 30009 24355 30067 24361
rect 30193 24327 30251 24333
rect 30193 24324 30205 24327
rect 28368 24296 30205 24324
rect 20901 24287 20959 24293
rect 30193 24293 30205 24296
rect 30239 24293 30251 24327
rect 30193 24287 30251 24293
rect 18874 24256 18880 24268
rect 16500 24228 17724 24256
rect 17788 24228 18880 24256
rect 16500 24200 16528 24228
rect 12526 24188 12532 24200
rect 12487 24160 12532 24188
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13078 24188 13084 24200
rect 13035 24160 13084 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13354 24188 13360 24200
rect 13315 24160 13360 24188
rect 13354 24148 13360 24160
rect 13412 24148 13418 24200
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 14783 24160 16037 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 16482 24188 16488 24200
rect 16347 24160 16488 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 13170 24120 13176 24132
rect 13131 24092 13176 24120
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 13265 24123 13323 24129
rect 13265 24089 13277 24123
rect 13311 24120 13323 24123
rect 13446 24120 13452 24132
rect 13311 24092 13452 24120
rect 13311 24089 13323 24092
rect 13265 24083 13323 24089
rect 13446 24080 13452 24092
rect 13504 24080 13510 24132
rect 16040 24120 16068 24151
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 16942 24148 16948 24200
rect 17000 24188 17006 24200
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17000 24160 17325 24188
rect 17000 24148 17006 24160
rect 17313 24157 17325 24160
rect 17359 24157 17371 24191
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17313 24151 17371 24157
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17696 24197 17724 24228
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 19334 24256 19340 24268
rect 19260 24228 19340 24256
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 16574 24120 16580 24132
rect 16040 24092 16580 24120
rect 16574 24080 16580 24092
rect 16632 24120 16638 24132
rect 17034 24120 17040 24132
rect 16632 24092 17040 24120
rect 16632 24080 16638 24092
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 17218 24080 17224 24132
rect 17276 24120 17282 24132
rect 17589 24123 17647 24129
rect 17589 24120 17601 24123
rect 17276 24092 17601 24120
rect 17276 24080 17282 24092
rect 17589 24089 17601 24092
rect 17635 24089 17647 24123
rect 17696 24120 17724 24151
rect 17770 24148 17776 24200
rect 17828 24188 17834 24200
rect 19260 24197 19288 24228
rect 19334 24216 19340 24228
rect 19392 24216 19398 24268
rect 21542 24256 21548 24268
rect 20548 24228 21548 24256
rect 18509 24191 18567 24197
rect 18509 24188 18521 24191
rect 17828 24160 18521 24188
rect 17828 24148 17834 24160
rect 18509 24157 18521 24160
rect 18555 24157 18567 24191
rect 18509 24151 18567 24157
rect 19245 24191 19303 24197
rect 19245 24157 19257 24191
rect 19291 24157 19303 24191
rect 19426 24188 19432 24200
rect 19387 24160 19432 24188
rect 19245 24151 19303 24157
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 19886 24188 19892 24200
rect 19847 24160 19892 24188
rect 19886 24148 19892 24160
rect 19944 24148 19950 24200
rect 20070 24188 20076 24200
rect 20031 24160 20076 24188
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20548 24197 20576 24228
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 21729 24259 21787 24265
rect 21729 24225 21741 24259
rect 21775 24256 21787 24259
rect 22186 24256 22192 24268
rect 21775 24228 22192 24256
rect 21775 24225 21787 24228
rect 21729 24219 21787 24225
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 22462 24216 22468 24268
rect 22520 24256 22526 24268
rect 23661 24259 23719 24265
rect 23661 24256 23673 24259
rect 22520 24228 23673 24256
rect 22520 24216 22526 24228
rect 23661 24225 23673 24228
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 30668 24265 30696 24364
rect 32766 24352 32772 24404
rect 32824 24392 32830 24404
rect 33505 24395 33563 24401
rect 33505 24392 33517 24395
rect 32824 24364 33517 24392
rect 32824 24352 32830 24364
rect 33505 24361 33517 24364
rect 33551 24392 33563 24395
rect 34698 24392 34704 24404
rect 33551 24364 34704 24392
rect 33551 24361 33563 24364
rect 33505 24355 33563 24361
rect 34698 24352 34704 24364
rect 34756 24352 34762 24404
rect 24489 24259 24547 24265
rect 24489 24256 24501 24259
rect 24176 24228 24501 24256
rect 24176 24216 24182 24228
rect 24489 24225 24501 24228
rect 24535 24225 24547 24259
rect 24489 24219 24547 24225
rect 30653 24259 30711 24265
rect 30653 24225 30665 24259
rect 30699 24256 30711 24259
rect 31202 24256 31208 24268
rect 30699 24228 31208 24256
rect 30699 24225 30711 24228
rect 30653 24219 30711 24225
rect 31202 24216 31208 24228
rect 31260 24216 31266 24268
rect 20538 24191 20596 24197
rect 20538 24157 20550 24191
rect 20584 24157 20596 24191
rect 20538 24151 20596 24157
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24188 20775 24191
rect 20806 24188 20812 24200
rect 20763 24160 20812 24188
rect 20763 24157 20775 24160
rect 20717 24151 20775 24157
rect 20806 24148 20812 24160
rect 20864 24148 20870 24200
rect 22002 24188 22008 24200
rect 21963 24160 22008 24188
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 24026 24188 24032 24200
rect 23523 24160 24032 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24188 24639 24191
rect 24670 24188 24676 24200
rect 24627 24160 24676 24188
rect 24627 24157 24639 24160
rect 24581 24151 24639 24157
rect 17696 24092 18552 24120
rect 17589 24083 17647 24089
rect 18524 24064 18552 24092
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 19904 24120 19932 24148
rect 19208 24092 19932 24120
rect 23569 24123 23627 24129
rect 19208 24080 19214 24092
rect 23569 24089 23581 24123
rect 23615 24120 23627 24123
rect 24596 24120 24624 24151
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24157 26295 24191
rect 27430 24188 27436 24200
rect 27391 24160 27436 24188
rect 26237 24151 26295 24157
rect 23615 24092 24624 24120
rect 25409 24123 25467 24129
rect 23615 24089 23627 24092
rect 23569 24083 23627 24089
rect 25409 24089 25421 24123
rect 25455 24120 25467 24123
rect 26050 24120 26056 24132
rect 25455 24092 26056 24120
rect 25455 24089 25467 24092
rect 25409 24083 25467 24089
rect 26050 24080 26056 24092
rect 26108 24080 26114 24132
rect 26252 24120 26280 24151
rect 27430 24148 27436 24160
rect 27488 24148 27494 24200
rect 27706 24197 27712 24200
rect 27700 24188 27712 24197
rect 27667 24160 27712 24188
rect 27700 24151 27712 24160
rect 27706 24148 27712 24151
rect 27764 24148 27770 24200
rect 29822 24188 29828 24200
rect 29783 24160 29828 24188
rect 29822 24148 29828 24160
rect 29880 24148 29886 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30926 24188 30932 24200
rect 30887 24160 30932 24188
rect 30009 24151 30067 24157
rect 28442 24120 28448 24132
rect 26252 24092 28448 24120
rect 28442 24080 28448 24092
rect 28500 24080 28506 24132
rect 30024 24120 30052 24151
rect 30926 24148 30932 24160
rect 30984 24148 30990 24200
rect 31662 24148 31668 24200
rect 31720 24188 31726 24200
rect 32125 24191 32183 24197
rect 32125 24188 32137 24191
rect 31720 24160 32137 24188
rect 31720 24148 31726 24160
rect 32125 24157 32137 24160
rect 32171 24188 32183 24191
rect 32171 24160 33088 24188
rect 32171 24157 32183 24160
rect 32125 24151 32183 24157
rect 33060 24132 33088 24160
rect 30834 24120 30840 24132
rect 30024 24092 30840 24120
rect 30834 24080 30840 24092
rect 30892 24120 30898 24132
rect 31294 24120 31300 24132
rect 30892 24092 31300 24120
rect 30892 24080 30898 24092
rect 31294 24080 31300 24092
rect 31352 24080 31358 24132
rect 32392 24123 32450 24129
rect 32392 24089 32404 24123
rect 32438 24120 32450 24123
rect 32950 24120 32956 24132
rect 32438 24092 32956 24120
rect 32438 24089 32450 24092
rect 32392 24083 32450 24089
rect 32950 24080 32956 24092
rect 33008 24080 33014 24132
rect 33042 24080 33048 24132
rect 33100 24080 33106 24132
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 12894 24012 12900 24064
rect 12952 24052 12958 24064
rect 13541 24055 13599 24061
rect 13541 24052 13553 24055
rect 12952 24024 13553 24052
rect 12952 24012 12958 24024
rect 13541 24021 13553 24024
rect 13587 24021 13599 24055
rect 13541 24015 13599 24021
rect 18230 24012 18236 24064
rect 18288 24052 18294 24064
rect 18325 24055 18383 24061
rect 18325 24052 18337 24055
rect 18288 24024 18337 24052
rect 18288 24012 18294 24024
rect 18325 24021 18337 24024
rect 18371 24021 18383 24055
rect 18325 24015 18383 24021
rect 18506 24012 18512 24064
rect 18564 24012 18570 24064
rect 19978 24052 19984 24064
rect 19939 24024 19984 24052
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20162 24012 20168 24064
rect 20220 24052 20226 24064
rect 23109 24055 23167 24061
rect 23109 24052 23121 24055
rect 20220 24024 23121 24052
rect 20220 24012 20226 24024
rect 23109 24021 23121 24024
rect 23155 24021 23167 24055
rect 23109 24015 23167 24021
rect 25590 24012 25596 24064
rect 25648 24061 25654 24064
rect 25648 24055 25667 24061
rect 25655 24021 25667 24055
rect 25774 24052 25780 24064
rect 25735 24024 25780 24052
rect 25648 24015 25667 24021
rect 25648 24012 25654 24015
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 27706 24012 27712 24064
rect 27764 24052 27770 24064
rect 27890 24052 27896 24064
rect 27764 24024 27896 24052
rect 27764 24012 27770 24024
rect 27890 24012 27896 24024
rect 27948 24012 27954 24064
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 28534 24052 28540 24064
rect 28408 24024 28540 24052
rect 28408 24012 28414 24024
rect 28534 24012 28540 24024
rect 28592 24052 28598 24064
rect 28813 24055 28871 24061
rect 28813 24052 28825 24055
rect 28592 24024 28825 24052
rect 28592 24012 28598 24024
rect 28813 24021 28825 24024
rect 28859 24021 28871 24055
rect 28813 24015 28871 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 13170 23808 13176 23860
rect 13228 23848 13234 23860
rect 13909 23851 13967 23857
rect 13909 23848 13921 23851
rect 13228 23820 13921 23848
rect 13228 23808 13234 23820
rect 13909 23817 13921 23820
rect 13955 23817 13967 23851
rect 13909 23811 13967 23817
rect 14277 23851 14335 23857
rect 14277 23817 14289 23851
rect 14323 23848 14335 23851
rect 15838 23848 15844 23860
rect 14323 23820 15844 23848
rect 14323 23817 14335 23820
rect 14277 23811 14335 23817
rect 12060 23783 12118 23789
rect 12060 23749 12072 23783
rect 12106 23780 12118 23783
rect 12342 23780 12348 23792
rect 12106 23752 12348 23780
rect 12106 23749 12118 23752
rect 12060 23743 12118 23749
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 11790 23712 11796 23724
rect 11751 23684 11796 23712
rect 11790 23672 11796 23684
rect 11848 23672 11854 23724
rect 13173 23579 13231 23585
rect 13173 23545 13185 23579
rect 13219 23576 13231 23579
rect 13446 23576 13452 23588
rect 13219 23548 13452 23576
rect 13219 23545 13231 23548
rect 13173 23539 13231 23545
rect 13446 23536 13452 23548
rect 13504 23576 13510 23588
rect 14292 23576 14320 23811
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17037 23851 17095 23857
rect 17037 23848 17049 23851
rect 16816 23820 17049 23848
rect 16816 23808 16822 23820
rect 17037 23817 17049 23820
rect 17083 23817 17095 23851
rect 17037 23811 17095 23817
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 21269 23851 21327 23857
rect 21269 23848 21281 23851
rect 18656 23820 21281 23848
rect 18656 23808 18662 23820
rect 21269 23817 21281 23820
rect 21315 23817 21327 23851
rect 21269 23811 21327 23817
rect 21910 23808 21916 23860
rect 21968 23848 21974 23860
rect 22021 23851 22079 23857
rect 22021 23848 22033 23851
rect 21968 23820 22033 23848
rect 21968 23808 21974 23820
rect 22021 23817 22033 23820
rect 22067 23817 22079 23851
rect 22021 23811 22079 23817
rect 24302 23808 24308 23860
rect 24360 23848 24366 23860
rect 24762 23848 24768 23860
rect 24360 23820 24768 23848
rect 24360 23808 24366 23820
rect 24762 23808 24768 23820
rect 24820 23848 24826 23860
rect 26973 23851 27031 23857
rect 24820 23820 26188 23848
rect 24820 23808 24826 23820
rect 19978 23780 19984 23792
rect 14568 23752 19984 23780
rect 14568 23653 14596 23752
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 20070 23740 20076 23792
rect 20128 23780 20134 23792
rect 20441 23783 20499 23789
rect 20441 23780 20453 23783
rect 20128 23752 20453 23780
rect 20128 23740 20134 23752
rect 20441 23749 20453 23752
rect 20487 23749 20499 23783
rect 20441 23743 20499 23749
rect 21821 23783 21879 23789
rect 21821 23749 21833 23783
rect 21867 23780 21879 23783
rect 21867 23752 21901 23780
rect 22066 23752 24348 23780
rect 21867 23749 21879 23752
rect 21821 23743 21879 23749
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23712 15347 23715
rect 15654 23712 15660 23724
rect 15335 23684 15660 23712
rect 15335 23681 15347 23684
rect 15289 23675 15347 23681
rect 15654 23672 15660 23684
rect 15712 23712 15718 23724
rect 16206 23712 16212 23724
rect 15712 23684 16212 23712
rect 15712 23672 15718 23684
rect 16206 23672 16212 23684
rect 16264 23672 16270 23724
rect 17862 23712 17868 23724
rect 17052 23684 17868 23712
rect 14369 23647 14427 23653
rect 14369 23613 14381 23647
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 15562 23644 15568 23656
rect 15523 23616 15568 23644
rect 14553 23607 14611 23613
rect 13504 23548 14320 23576
rect 14384 23576 14412 23607
rect 15562 23604 15568 23616
rect 15620 23644 15626 23656
rect 16942 23644 16948 23656
rect 15620 23616 16948 23644
rect 15620 23604 15626 23616
rect 16942 23604 16948 23616
rect 17000 23644 17006 23656
rect 17052 23644 17080 23684
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 18046 23712 18052 23724
rect 18007 23684 18052 23712
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 18138 23672 18144 23724
rect 18196 23712 18202 23724
rect 18279 23715 18337 23721
rect 18196 23684 18241 23712
rect 18196 23672 18202 23684
rect 18279 23681 18291 23715
rect 18325 23712 18337 23715
rect 18506 23712 18512 23724
rect 18325 23684 18512 23712
rect 18325 23681 18337 23684
rect 18279 23675 18337 23681
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 20088 23712 20116 23740
rect 19475 23684 20116 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 20162 23672 20168 23724
rect 20220 23712 20226 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20220 23684 20269 23712
rect 20220 23672 20226 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20438 23712 20444 23714
rect 20257 23675 20315 23681
rect 20364 23684 20444 23712
rect 17000 23616 17080 23644
rect 17129 23647 17187 23653
rect 17000 23604 17006 23616
rect 17129 23613 17141 23647
rect 17175 23613 17187 23647
rect 17129 23607 17187 23613
rect 17313 23647 17371 23653
rect 17313 23613 17325 23647
rect 17359 23644 17371 23647
rect 18414 23644 18420 23656
rect 17359 23616 18420 23644
rect 17359 23613 17371 23616
rect 17313 23607 17371 23613
rect 14642 23576 14648 23588
rect 14384 23548 14648 23576
rect 13504 23536 13510 23548
rect 14642 23536 14648 23548
rect 14700 23576 14706 23588
rect 17144 23576 17172 23607
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 20036 23616 20085 23644
rect 20036 23604 20042 23616
rect 20073 23613 20085 23616
rect 20119 23644 20131 23647
rect 20364 23644 20392 23684
rect 20438 23662 20444 23684
rect 20496 23662 20502 23714
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 20901 23715 20959 23721
rect 20901 23712 20913 23715
rect 20772 23684 20913 23712
rect 20772 23672 20778 23684
rect 20901 23681 20913 23684
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21266 23712 21272 23724
rect 21131 23684 21272 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 21836 23712 21864 23743
rect 22066 23712 22094 23752
rect 21784 23684 22094 23712
rect 21784 23672 21790 23684
rect 22186 23672 22192 23724
rect 22244 23712 22250 23724
rect 22649 23715 22707 23721
rect 22649 23712 22661 23715
rect 22244 23684 22661 23712
rect 22244 23672 22250 23684
rect 22649 23681 22661 23684
rect 22695 23681 22707 23715
rect 22830 23712 22836 23724
rect 22791 23684 22836 23712
rect 22649 23675 22707 23681
rect 22830 23672 22836 23684
rect 22888 23712 22894 23724
rect 24320 23721 24348 23752
rect 25314 23740 25320 23792
rect 25372 23780 25378 23792
rect 25682 23780 25688 23792
rect 25372 23752 25688 23780
rect 25372 23740 25378 23752
rect 25682 23740 25688 23752
rect 25740 23740 25746 23792
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 22888 23684 23673 23712
rect 22888 23672 22894 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 24305 23715 24363 23721
rect 24305 23681 24317 23715
rect 24351 23681 24363 23715
rect 24305 23675 24363 23681
rect 25225 23715 25283 23721
rect 25225 23681 25237 23715
rect 25271 23712 25283 23715
rect 25332 23712 25360 23740
rect 25271 23684 25360 23712
rect 25409 23715 25467 23721
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 25409 23681 25421 23715
rect 25455 23712 25467 23715
rect 25498 23712 25504 23724
rect 25455 23684 25504 23712
rect 25455 23681 25467 23684
rect 25409 23675 25467 23681
rect 20119 23616 20392 23644
rect 20119 23613 20131 23616
rect 20073 23607 20131 23613
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22741 23647 22799 23653
rect 22741 23644 22753 23647
rect 21968 23616 22753 23644
rect 21968 23604 21974 23616
rect 22741 23613 22753 23616
rect 22787 23613 22799 23647
rect 23676 23644 23704 23675
rect 25498 23672 25504 23684
rect 25556 23672 25562 23724
rect 25958 23712 25964 23724
rect 25919 23684 25964 23712
rect 25958 23672 25964 23684
rect 26016 23672 26022 23724
rect 26160 23721 26188 23820
rect 26973 23817 26985 23851
rect 27019 23848 27031 23851
rect 27982 23848 27988 23860
rect 27019 23820 27988 23848
rect 27019 23817 27031 23820
rect 26973 23811 27031 23817
rect 27982 23808 27988 23820
rect 28040 23848 28046 23860
rect 28077 23851 28135 23857
rect 28077 23848 28089 23851
rect 28040 23820 28089 23848
rect 28040 23808 28046 23820
rect 28077 23817 28089 23820
rect 28123 23817 28135 23851
rect 28077 23811 28135 23817
rect 28626 23808 28632 23860
rect 28684 23848 28690 23860
rect 28684 23820 31984 23848
rect 28684 23808 28690 23820
rect 27341 23783 27399 23789
rect 27341 23780 27353 23783
rect 26252 23752 27353 23780
rect 26145 23715 26203 23721
rect 26145 23681 26157 23715
rect 26191 23681 26203 23715
rect 26145 23675 26203 23681
rect 23676 23616 23980 23644
rect 22741 23607 22799 23613
rect 14700 23548 17172 23576
rect 14700 23536 14706 23548
rect 20438 23536 20444 23588
rect 20496 23576 20502 23588
rect 22189 23579 22247 23585
rect 22189 23576 22201 23579
rect 20496 23548 22201 23576
rect 20496 23536 20502 23548
rect 22189 23545 22201 23548
rect 22235 23545 22247 23579
rect 23842 23576 23848 23588
rect 23803 23548 23848 23576
rect 22189 23539 22247 23545
rect 23842 23536 23848 23548
rect 23900 23536 23906 23588
rect 23952 23576 23980 23616
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 25096 23616 25145 23644
rect 25096 23604 25102 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25317 23647 25375 23653
rect 25317 23644 25329 23647
rect 25133 23607 25191 23613
rect 25240 23616 25329 23644
rect 25240 23588 25268 23616
rect 25317 23613 25329 23616
rect 25363 23644 25375 23647
rect 26252 23644 26280 23752
rect 27341 23749 27353 23752
rect 27387 23749 27399 23783
rect 27341 23743 27399 23749
rect 28994 23740 29000 23792
rect 29052 23780 29058 23792
rect 29914 23780 29920 23792
rect 29052 23752 29920 23780
rect 29052 23740 29058 23752
rect 29914 23740 29920 23752
rect 29972 23780 29978 23792
rect 30558 23780 30564 23792
rect 29972 23752 30564 23780
rect 29972 23740 29978 23752
rect 30558 23740 30564 23752
rect 30616 23740 30622 23792
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23681 27491 23715
rect 27433 23675 27491 23681
rect 28074 23715 28132 23721
rect 28074 23681 28086 23715
rect 28120 23712 28132 23715
rect 28166 23712 28172 23724
rect 28120 23684 28172 23712
rect 28120 23681 28132 23684
rect 28074 23675 28132 23681
rect 25363 23616 26280 23644
rect 25363 23613 25375 23616
rect 25317 23607 25375 23613
rect 23952 23548 25084 23576
rect 16666 23508 16672 23520
rect 16627 23480 16672 23508
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 18417 23511 18475 23517
rect 18417 23508 18429 23511
rect 17000 23480 18429 23508
rect 17000 23468 17006 23480
rect 18417 23477 18429 23480
rect 18463 23477 18475 23511
rect 19518 23508 19524 23520
rect 19479 23480 19524 23508
rect 18417 23471 18475 23477
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 21085 23511 21143 23517
rect 21085 23508 21097 23511
rect 21048 23480 21097 23508
rect 21048 23468 21054 23480
rect 21085 23477 21097 23480
rect 21131 23508 21143 23511
rect 21818 23508 21824 23520
rect 21131 23480 21824 23508
rect 21131 23477 21143 23480
rect 21085 23471 21143 23477
rect 21818 23468 21824 23480
rect 21876 23468 21882 23520
rect 22005 23511 22063 23517
rect 22005 23477 22017 23511
rect 22051 23508 22063 23511
rect 22554 23508 22560 23520
rect 22051 23480 22560 23508
rect 22051 23477 22063 23480
rect 22005 23471 22063 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 24302 23468 24308 23520
rect 24360 23508 24366 23520
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24360 23480 24409 23508
rect 24360 23468 24366 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 24762 23468 24768 23520
rect 24820 23508 24826 23520
rect 24949 23511 25007 23517
rect 24949 23508 24961 23511
rect 24820 23480 24961 23508
rect 24820 23468 24826 23480
rect 24949 23477 24961 23480
rect 24995 23477 25007 23511
rect 25056 23508 25084 23548
rect 25222 23536 25228 23588
rect 25280 23536 25286 23588
rect 27172 23576 27200 23675
rect 27448 23644 27476 23675
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 29181 23715 29239 23721
rect 29181 23681 29193 23715
rect 29227 23681 29239 23715
rect 29181 23675 29239 23681
rect 28350 23644 28356 23656
rect 27448 23616 28356 23644
rect 28350 23604 28356 23616
rect 28408 23604 28414 23656
rect 28534 23644 28540 23656
rect 28495 23616 28540 23644
rect 28534 23604 28540 23616
rect 28592 23644 28598 23656
rect 29196 23644 29224 23675
rect 29270 23672 29276 23724
rect 29328 23712 29334 23724
rect 30285 23715 30343 23721
rect 29328 23684 29373 23712
rect 29328 23672 29334 23684
rect 30285 23681 30297 23715
rect 30331 23712 30343 23715
rect 31754 23712 31760 23724
rect 30331 23684 31760 23712
rect 30331 23681 30343 23684
rect 30285 23675 30343 23681
rect 28592 23616 29224 23644
rect 28592 23604 28598 23616
rect 28445 23579 28503 23585
rect 28445 23576 28457 23579
rect 27172 23548 28457 23576
rect 28445 23545 28457 23548
rect 28491 23576 28503 23579
rect 28810 23576 28816 23588
rect 28491 23548 28816 23576
rect 28491 23545 28503 23548
rect 28445 23539 28503 23545
rect 28810 23536 28816 23548
rect 28868 23576 28874 23588
rect 30300 23576 30328 23675
rect 31754 23672 31760 23684
rect 31812 23672 31818 23724
rect 30558 23644 30564 23656
rect 30471 23616 30564 23644
rect 30558 23604 30564 23616
rect 30616 23604 30622 23656
rect 31956 23644 31984 23820
rect 32950 23808 32956 23860
rect 33008 23848 33014 23860
rect 33321 23851 33379 23857
rect 33321 23848 33333 23851
rect 33008 23820 33333 23848
rect 33008 23808 33014 23820
rect 33321 23817 33333 23820
rect 33367 23817 33379 23851
rect 33321 23811 33379 23817
rect 33410 23808 33416 23860
rect 33468 23848 33474 23860
rect 33468 23820 34100 23848
rect 33468 23808 33474 23820
rect 32030 23740 32036 23792
rect 32088 23780 32094 23792
rect 32490 23780 32496 23792
rect 32088 23752 32352 23780
rect 32088 23740 32094 23752
rect 32122 23712 32128 23724
rect 32083 23684 32128 23712
rect 32122 23672 32128 23684
rect 32180 23672 32186 23724
rect 32324 23721 32352 23752
rect 32416 23752 32496 23780
rect 32416 23721 32444 23752
rect 32490 23740 32496 23752
rect 32548 23740 32554 23792
rect 32861 23783 32919 23789
rect 32861 23749 32873 23783
rect 32907 23780 32919 23783
rect 32907 23752 33732 23780
rect 32907 23749 32919 23752
rect 32861 23743 32919 23749
rect 32309 23715 32367 23721
rect 32309 23681 32321 23715
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 32401 23715 32459 23721
rect 32401 23681 32413 23715
rect 32447 23681 32459 23715
rect 32401 23675 32459 23681
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23714 32735 23715
rect 32766 23714 32772 23724
rect 32723 23686 32772 23714
rect 32723 23681 32735 23686
rect 32677 23675 32735 23681
rect 32766 23672 32772 23686
rect 32824 23672 32830 23724
rect 32950 23672 32956 23724
rect 33008 23712 33014 23724
rect 33704 23721 33732 23752
rect 33597 23715 33655 23721
rect 33597 23712 33609 23715
rect 33008 23684 33609 23712
rect 33008 23672 33014 23684
rect 33597 23681 33609 23684
rect 33643 23681 33655 23715
rect 33597 23675 33655 23681
rect 33689 23715 33747 23721
rect 33689 23681 33701 23715
rect 33735 23681 33747 23715
rect 33689 23675 33747 23681
rect 33778 23672 33784 23724
rect 33836 23712 33842 23724
rect 33941 23715 33999 23721
rect 33836 23684 33881 23712
rect 33836 23672 33842 23684
rect 33941 23681 33953 23715
rect 33987 23712 33999 23715
rect 34072 23712 34100 23820
rect 34422 23712 34428 23724
rect 33987 23684 34100 23712
rect 34383 23684 34428 23712
rect 33987 23681 33999 23684
rect 33941 23675 33999 23681
rect 34422 23672 34428 23684
rect 34480 23672 34486 23724
rect 34609 23715 34667 23721
rect 34609 23681 34621 23715
rect 34655 23681 34667 23715
rect 34609 23675 34667 23681
rect 32493 23647 32551 23653
rect 32493 23644 32505 23647
rect 31956 23616 32505 23644
rect 32493 23613 32505 23616
rect 32539 23644 32551 23647
rect 32539 23616 34100 23644
rect 32539 23613 32551 23616
rect 32493 23607 32551 23613
rect 28868 23548 30328 23576
rect 30576 23576 30604 23604
rect 32766 23576 32772 23588
rect 30576 23548 32772 23576
rect 28868 23536 28874 23548
rect 32766 23536 32772 23548
rect 32824 23536 32830 23588
rect 32858 23536 32864 23588
rect 32916 23576 32922 23588
rect 33778 23576 33784 23588
rect 32916 23548 33784 23576
rect 32916 23536 32922 23548
rect 33778 23536 33784 23548
rect 33836 23536 33842 23588
rect 34072 23576 34100 23616
rect 34146 23604 34152 23656
rect 34204 23644 34210 23656
rect 34624 23644 34652 23675
rect 34204 23616 34652 23644
rect 34204 23604 34210 23616
rect 34422 23576 34428 23588
rect 34072 23548 34428 23576
rect 34422 23536 34428 23548
rect 34480 23536 34486 23588
rect 25961 23511 26019 23517
rect 25961 23508 25973 23511
rect 25056 23480 25973 23508
rect 24949 23471 25007 23477
rect 25961 23477 25973 23480
rect 26007 23477 26019 23511
rect 25961 23471 26019 23477
rect 27893 23511 27951 23517
rect 27893 23477 27905 23511
rect 27939 23508 27951 23511
rect 28258 23508 28264 23520
rect 27939 23480 28264 23508
rect 27939 23477 27951 23480
rect 27893 23471 27951 23477
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 28997 23511 29055 23517
rect 28997 23477 29009 23511
rect 29043 23508 29055 23511
rect 31386 23508 31392 23520
rect 29043 23480 31392 23508
rect 29043 23477 29055 23480
rect 28997 23471 29055 23477
rect 31386 23468 31392 23480
rect 31444 23468 31450 23520
rect 32122 23468 32128 23520
rect 32180 23508 32186 23520
rect 34517 23511 34575 23517
rect 34517 23508 34529 23511
rect 32180 23480 34529 23508
rect 32180 23468 32186 23480
rect 34517 23477 34529 23480
rect 34563 23477 34575 23511
rect 34517 23471 34575 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 16666 23304 16672 23316
rect 13648 23276 16672 23304
rect 13541 23239 13599 23245
rect 13541 23236 13553 23239
rect 11532 23208 13553 23236
rect 11532 23109 11560 23208
rect 13541 23205 13553 23208
rect 13587 23205 13599 23239
rect 13541 23199 13599 23205
rect 12161 23171 12219 23177
rect 12161 23137 12173 23171
rect 12207 23168 12219 23171
rect 12434 23168 12440 23180
rect 12207 23140 12440 23168
rect 12207 23137 12219 23140
rect 12161 23131 12219 23137
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23069 11483 23103
rect 11425 23063 11483 23069
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 11440 23032 11468 23063
rect 12176 23032 12204 23131
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 13648 23168 13676 23276
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 17681 23307 17739 23313
rect 17681 23273 17693 23307
rect 17727 23304 17739 23307
rect 18046 23304 18052 23316
rect 17727 23276 18052 23304
rect 17727 23273 17739 23276
rect 17681 23267 17739 23273
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 19610 23304 19616 23316
rect 18156 23276 19616 23304
rect 15654 23236 15660 23248
rect 13188 23140 13676 23168
rect 14660 23208 15660 23236
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23100 12403 23103
rect 12894 23100 12900 23112
rect 12391 23072 12900 23100
rect 12391 23069 12403 23072
rect 12345 23063 12403 23069
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13078 23100 13084 23112
rect 13035 23072 13084 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 13188 23109 13216 23140
rect 13173 23103 13231 23109
rect 13173 23069 13185 23103
rect 13219 23069 13231 23103
rect 13354 23100 13360 23112
rect 13315 23072 13360 23100
rect 13173 23063 13231 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 14660 23109 14688 23208
rect 15654 23196 15660 23208
rect 15712 23196 15718 23248
rect 16574 23196 16580 23248
rect 16632 23236 16638 23248
rect 18156 23236 18184 23276
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 20438 23304 20444 23316
rect 20399 23276 20444 23304
rect 20438 23264 20444 23276
rect 20496 23264 20502 23316
rect 22922 23304 22928 23316
rect 22883 23276 22928 23304
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 24596 23276 25912 23304
rect 24596 23236 24624 23276
rect 16632 23208 18184 23236
rect 19260 23208 24624 23236
rect 25884 23236 25912 23276
rect 26142 23264 26148 23316
rect 26200 23304 26206 23316
rect 26329 23307 26387 23313
rect 26329 23304 26341 23307
rect 26200 23276 26341 23304
rect 26200 23264 26206 23276
rect 26329 23273 26341 23276
rect 26375 23273 26387 23307
rect 26329 23267 26387 23273
rect 30466 23264 30472 23316
rect 30524 23304 30530 23316
rect 30653 23307 30711 23313
rect 30653 23304 30665 23307
rect 30524 23276 30665 23304
rect 30524 23264 30530 23276
rect 30653 23273 30665 23276
rect 30699 23273 30711 23307
rect 34790 23304 34796 23316
rect 34751 23276 34796 23304
rect 30653 23267 30711 23273
rect 34790 23264 34796 23276
rect 34848 23264 34854 23316
rect 27062 23236 27068 23248
rect 25884 23208 27068 23236
rect 16632 23196 16638 23208
rect 14826 23128 14832 23180
rect 14884 23168 14890 23180
rect 16206 23168 16212 23180
rect 14884 23140 16212 23168
rect 14884 23128 14890 23140
rect 16206 23128 16212 23140
rect 16264 23168 16270 23180
rect 16945 23171 17003 23177
rect 16945 23168 16957 23171
rect 16264 23140 16957 23168
rect 16264 23128 16270 23140
rect 16945 23137 16957 23140
rect 16991 23168 17003 23171
rect 17034 23168 17040 23180
rect 16991 23140 17040 23168
rect 16991 23137 17003 23140
rect 16945 23131 17003 23137
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23168 17187 23171
rect 18046 23168 18052 23180
rect 17175 23140 18052 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 18046 23128 18052 23140
rect 18104 23128 18110 23180
rect 18322 23168 18328 23180
rect 18283 23140 18328 23168
rect 18322 23128 18328 23140
rect 18380 23128 18386 23180
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 14921 23103 14979 23109
rect 14921 23069 14933 23103
rect 14967 23069 14979 23103
rect 17052 23100 17080 23128
rect 17586 23100 17592 23112
rect 17052 23072 17592 23100
rect 14921 23063 14979 23069
rect 11440 23004 12204 23032
rect 13096 23032 13124 23060
rect 13265 23035 13323 23041
rect 13096 23004 13216 23032
rect 13188 22976 13216 23004
rect 13265 23001 13277 23035
rect 13311 23032 13323 23035
rect 13446 23032 13452 23044
rect 13311 23004 13452 23032
rect 13311 23001 13323 23004
rect 13265 22995 13323 23001
rect 13446 22992 13452 23004
rect 13504 22992 13510 23044
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22964 11759 22967
rect 13078 22964 13084 22976
rect 11747 22936 13084 22964
rect 11747 22933 11759 22936
rect 11701 22927 11759 22933
rect 13078 22924 13084 22936
rect 13136 22924 13142 22976
rect 13170 22924 13176 22976
rect 13228 22964 13234 22976
rect 14936 22964 14964 23063
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 18138 23060 18144 23112
rect 18196 23060 18202 23112
rect 19260 23109 19288 23208
rect 27062 23196 27068 23208
rect 27120 23196 27126 23248
rect 27522 23236 27528 23248
rect 27483 23208 27528 23236
rect 27522 23196 27528 23208
rect 27580 23196 27586 23248
rect 30374 23196 30380 23248
rect 30432 23236 30438 23248
rect 31113 23239 31171 23245
rect 31113 23236 31125 23239
rect 30432 23208 31125 23236
rect 30432 23196 30438 23208
rect 31113 23205 31125 23208
rect 31159 23205 31171 23239
rect 31113 23199 31171 23205
rect 19426 23128 19432 23180
rect 19484 23168 19490 23180
rect 19484 23140 19932 23168
rect 19484 23128 19490 23140
rect 19904 23112 19932 23140
rect 20162 23128 20168 23180
rect 20220 23168 20226 23180
rect 20441 23171 20499 23177
rect 20441 23168 20453 23171
rect 20220 23140 20453 23168
rect 20220 23128 20226 23140
rect 20441 23137 20453 23140
rect 20487 23137 20499 23171
rect 20441 23131 20499 23137
rect 20714 23128 20720 23180
rect 20772 23168 20778 23180
rect 21174 23168 21180 23180
rect 20772 23140 21180 23168
rect 20772 23128 20778 23140
rect 21174 23128 21180 23140
rect 21232 23168 21238 23180
rect 21913 23171 21971 23177
rect 21913 23168 21925 23171
rect 21232 23140 21925 23168
rect 21232 23128 21238 23140
rect 21913 23137 21925 23140
rect 21959 23137 21971 23171
rect 23750 23168 23756 23180
rect 21913 23131 21971 23137
rect 22940 23140 23756 23168
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19392 23072 19533 23100
rect 19392 23060 19398 23072
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 18049 23035 18107 23041
rect 18049 23001 18061 23035
rect 18095 23032 18107 23035
rect 18156 23032 18184 23060
rect 18598 23032 18604 23044
rect 18095 23004 18604 23032
rect 18095 23001 18107 23004
rect 18049 22995 18107 23001
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 19536 23032 19564 23063
rect 19610 23060 19616 23112
rect 19668 23100 19674 23112
rect 19668 23072 19713 23100
rect 19668 23060 19674 23072
rect 19886 23060 19892 23112
rect 19944 23100 19950 23112
rect 20349 23103 20407 23109
rect 20349 23100 20361 23103
rect 19944 23072 20361 23100
rect 19944 23060 19950 23072
rect 20349 23069 20361 23072
rect 20395 23069 20407 23103
rect 20622 23100 20628 23112
rect 20583 23072 20628 23100
rect 20349 23063 20407 23069
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 21637 23103 21695 23109
rect 21637 23069 21649 23103
rect 21683 23100 21695 23103
rect 21818 23100 21824 23112
rect 21683 23072 21824 23100
rect 21683 23069 21695 23072
rect 21637 23063 21695 23069
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 22940 23109 22968 23140
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 23845 23171 23903 23177
rect 23845 23137 23857 23171
rect 23891 23168 23903 23171
rect 24026 23168 24032 23180
rect 23891 23140 24032 23168
rect 23891 23137 23903 23140
rect 23845 23131 23903 23137
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 24762 23128 24768 23180
rect 24820 23168 24826 23180
rect 24820 23140 25084 23168
rect 24820 23128 24826 23140
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23100 23167 23103
rect 23198 23100 23204 23112
rect 23155 23072 23204 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 23584 23072 23888 23100
rect 23584 23032 23612 23072
rect 19536 23004 23612 23032
rect 23661 23035 23719 23041
rect 23661 23001 23673 23035
rect 23707 23032 23719 23035
rect 23750 23032 23756 23044
rect 23707 23004 23756 23032
rect 23707 23001 23719 23004
rect 23661 22995 23719 23001
rect 13228 22936 14964 22964
rect 16485 22967 16543 22973
rect 13228 22924 13234 22936
rect 16485 22933 16497 22967
rect 16531 22964 16543 22967
rect 16758 22964 16764 22976
rect 16531 22936 16764 22964
rect 16531 22933 16543 22936
rect 16485 22927 16543 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 16853 22967 16911 22973
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 17310 22964 17316 22976
rect 16899 22936 17316 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 17310 22924 17316 22936
rect 17368 22924 17374 22976
rect 17586 22924 17592 22976
rect 17644 22964 17650 22976
rect 18141 22967 18199 22973
rect 18141 22964 18153 22967
rect 17644 22936 18153 22964
rect 17644 22924 17650 22936
rect 18141 22933 18153 22936
rect 18187 22933 18199 22967
rect 18141 22927 18199 22933
rect 18322 22924 18328 22976
rect 18380 22964 18386 22976
rect 20809 22967 20867 22973
rect 20809 22964 20821 22967
rect 18380 22936 20821 22964
rect 18380 22924 18386 22936
rect 20809 22933 20821 22936
rect 20855 22933 20867 22967
rect 20809 22927 20867 22933
rect 22370 22924 22376 22976
rect 22428 22964 22434 22976
rect 23566 22964 23572 22976
rect 22428 22936 23572 22964
rect 22428 22924 22434 22936
rect 23566 22924 23572 22936
rect 23624 22964 23630 22976
rect 23676 22964 23704 22995
rect 23750 22992 23756 23004
rect 23808 22992 23814 23044
rect 23860 23032 23888 23072
rect 24854 23060 24860 23112
rect 24912 23100 24918 23112
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 24912 23072 24961 23100
rect 24912 23060 24918 23072
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 25056 23100 25084 23140
rect 29730 23128 29736 23180
rect 29788 23168 29794 23180
rect 30193 23171 30251 23177
rect 30193 23168 30205 23171
rect 29788 23140 30205 23168
rect 29788 23128 29794 23140
rect 30193 23137 30205 23140
rect 30239 23137 30251 23171
rect 31018 23168 31024 23180
rect 30193 23131 30251 23137
rect 30300 23140 31024 23168
rect 25205 23103 25263 23109
rect 25205 23100 25217 23103
rect 25056 23072 25217 23100
rect 24949 23063 25007 23069
rect 25205 23069 25217 23072
rect 25251 23069 25263 23103
rect 25205 23063 25263 23069
rect 25590 23060 25596 23112
rect 25648 23100 25654 23112
rect 29917 23103 29975 23109
rect 29917 23100 29929 23103
rect 25648 23072 29929 23100
rect 25648 23060 25654 23072
rect 29917 23069 29929 23072
rect 29963 23100 29975 23103
rect 30006 23100 30012 23112
rect 29963 23072 30012 23100
rect 29963 23069 29975 23072
rect 29917 23063 29975 23069
rect 30006 23060 30012 23072
rect 30064 23060 30070 23112
rect 30300 23109 30328 23140
rect 31018 23128 31024 23140
rect 31076 23168 31082 23180
rect 32490 23168 32496 23180
rect 31076 23140 32496 23168
rect 31076 23128 31082 23140
rect 32490 23128 32496 23140
rect 32548 23128 32554 23180
rect 32950 23168 32956 23180
rect 32692 23140 32956 23168
rect 30101 23103 30159 23109
rect 30101 23069 30113 23103
rect 30147 23069 30159 23103
rect 30101 23063 30159 23069
rect 30285 23103 30343 23109
rect 30285 23069 30297 23103
rect 30331 23069 30343 23103
rect 30285 23063 30343 23069
rect 27154 23032 27160 23044
rect 23860 23004 26188 23032
rect 27115 23004 27160 23032
rect 23624 22936 23704 22964
rect 23624 22924 23630 22936
rect 23842 22924 23848 22976
rect 23900 22964 23906 22976
rect 26050 22964 26056 22976
rect 23900 22936 26056 22964
rect 23900 22924 23906 22936
rect 26050 22924 26056 22936
rect 26108 22924 26114 22976
rect 26160 22964 26188 23004
rect 27154 22992 27160 23004
rect 27212 22992 27218 23044
rect 27522 22992 27528 23044
rect 27580 23032 27586 23044
rect 28445 23035 28503 23041
rect 28445 23032 28457 23035
rect 27580 23004 28457 23032
rect 27580 22992 27586 23004
rect 28445 23001 28457 23004
rect 28491 23001 28503 23035
rect 28626 23032 28632 23044
rect 28587 23004 28632 23032
rect 28445 22995 28503 23001
rect 28626 22992 28632 23004
rect 28684 22992 28690 23044
rect 30116 23032 30144 23063
rect 30466 23060 30472 23112
rect 30524 23100 30530 23112
rect 30926 23100 30932 23112
rect 30524 23072 30932 23100
rect 30524 23060 30530 23072
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 31386 23100 31392 23112
rect 31347 23072 31392 23100
rect 31386 23060 31392 23072
rect 31444 23060 31450 23112
rect 32122 23100 32128 23112
rect 31726 23072 32128 23100
rect 30374 23032 30380 23044
rect 30116 23004 30380 23032
rect 30374 22992 30380 23004
rect 30432 22992 30438 23044
rect 30558 22992 30564 23044
rect 30616 23032 30622 23044
rect 31113 23035 31171 23041
rect 31113 23032 31125 23035
rect 30616 23004 31125 23032
rect 30616 22992 30622 23004
rect 31113 23001 31125 23004
rect 31159 23001 31171 23035
rect 31113 22995 31171 23001
rect 31202 22992 31208 23044
rect 31260 23032 31266 23044
rect 31726 23032 31754 23072
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 32306 23100 32312 23112
rect 32267 23072 32312 23100
rect 32306 23060 32312 23072
rect 32364 23060 32370 23112
rect 32398 23060 32404 23112
rect 32456 23100 32462 23112
rect 32692 23109 32720 23140
rect 32950 23128 32956 23140
rect 33008 23168 33014 23180
rect 33597 23171 33655 23177
rect 33597 23168 33609 23171
rect 33008 23140 33609 23168
rect 33008 23128 33014 23140
rect 33597 23137 33609 23140
rect 33643 23137 33655 23171
rect 33597 23131 33655 23137
rect 32677 23103 32735 23109
rect 32456 23072 32501 23100
rect 32456 23060 32462 23072
rect 32677 23069 32689 23103
rect 32723 23069 32735 23103
rect 33318 23100 33324 23112
rect 33279 23072 33324 23100
rect 32677 23063 32735 23069
rect 33318 23060 33324 23072
rect 33376 23060 33382 23112
rect 34698 23100 34704 23112
rect 34659 23072 34704 23100
rect 34698 23060 34704 23072
rect 34756 23060 34762 23112
rect 31260 23004 31754 23032
rect 31260 22992 31266 23004
rect 27617 22967 27675 22973
rect 27617 22964 27629 22967
rect 26160 22936 27629 22964
rect 27617 22933 27629 22936
rect 27663 22933 27675 22967
rect 27617 22927 27675 22933
rect 28813 22967 28871 22973
rect 28813 22933 28825 22967
rect 28859 22964 28871 22967
rect 29638 22964 29644 22976
rect 28859 22936 29644 22964
rect 28859 22933 28871 22936
rect 28813 22927 28871 22933
rect 29638 22924 29644 22936
rect 29696 22924 29702 22976
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 31297 22967 31355 22973
rect 31297 22964 31309 22967
rect 30156 22936 31309 22964
rect 30156 22924 30162 22936
rect 31297 22933 31309 22936
rect 31343 22933 31355 22967
rect 32858 22964 32864 22976
rect 32819 22936 32864 22964
rect 31297 22927 31355 22933
rect 32858 22924 32864 22936
rect 32916 22924 32922 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 14826 22760 14832 22772
rect 14787 22732 14832 22760
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 18322 22760 18328 22772
rect 15580 22732 18328 22760
rect 12802 22692 12808 22704
rect 11992 22664 12808 22692
rect 11790 22584 11796 22636
rect 11848 22624 11854 22636
rect 11992 22633 12020 22664
rect 12802 22652 12808 22664
rect 12860 22652 12866 22704
rect 13078 22652 13084 22704
rect 13136 22692 13142 22704
rect 13136 22664 14044 22692
rect 13136 22652 13142 22664
rect 14016 22633 14044 22664
rect 11977 22627 12035 22633
rect 11977 22624 11989 22627
rect 11848 22596 11989 22624
rect 11848 22584 11854 22596
rect 11977 22593 11989 22596
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 12244 22627 12302 22633
rect 12244 22593 12256 22627
rect 12290 22624 12302 22627
rect 14001 22627 14059 22633
rect 12290 22596 13860 22624
rect 12290 22593 12302 22596
rect 12244 22587 12302 22593
rect 13832 22497 13860 22596
rect 14001 22593 14013 22627
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 14274 22516 14280 22568
rect 14332 22556 14338 22568
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14332 22528 14933 22556
rect 14332 22516 14338 22528
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 15105 22559 15163 22565
rect 15105 22525 15117 22559
rect 15151 22556 15163 22559
rect 15580 22556 15608 22732
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 21082 22760 21088 22772
rect 19444 22732 21088 22760
rect 15654 22652 15660 22704
rect 15712 22692 15718 22704
rect 17488 22695 17546 22701
rect 15712 22664 17356 22692
rect 15712 22652 15718 22664
rect 15746 22624 15752 22636
rect 15707 22596 15752 22624
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 15151 22528 15608 22556
rect 15856 22556 15884 22587
rect 16298 22584 16304 22636
rect 16356 22624 16362 22636
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 16356 22596 17233 22624
rect 16356 22584 16362 22596
rect 17221 22593 17233 22596
rect 17267 22593 17279 22627
rect 17328 22624 17356 22664
rect 17488 22661 17500 22695
rect 17534 22692 17546 22695
rect 18230 22692 18236 22704
rect 17534 22664 18236 22692
rect 17534 22661 17546 22664
rect 17488 22655 17546 22661
rect 18230 22652 18236 22664
rect 18288 22652 18294 22704
rect 19242 22692 19248 22704
rect 18340 22664 19248 22692
rect 18340 22624 18368 22664
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 19334 22624 19340 22636
rect 17328 22596 18368 22624
rect 19295 22596 19340 22624
rect 17221 22587 17279 22593
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 17126 22556 17132 22568
rect 15856 22528 17132 22556
rect 15151 22525 15163 22528
rect 15105 22519 15163 22525
rect 17126 22516 17132 22528
rect 17184 22516 17190 22568
rect 13817 22491 13875 22497
rect 13817 22457 13829 22491
rect 13863 22457 13875 22491
rect 16666 22488 16672 22500
rect 13817 22451 13875 22457
rect 14292 22460 16672 22488
rect 13357 22423 13415 22429
rect 13357 22389 13369 22423
rect 13403 22420 13415 22423
rect 13446 22420 13452 22432
rect 13403 22392 13452 22420
rect 13403 22389 13415 22392
rect 13357 22383 13415 22389
rect 13446 22380 13452 22392
rect 13504 22420 13510 22432
rect 14292 22420 14320 22460
rect 16666 22448 16672 22460
rect 16724 22448 16730 22500
rect 14458 22420 14464 22432
rect 13504 22392 14320 22420
rect 14419 22392 14464 22420
rect 13504 22380 13510 22392
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 16025 22423 16083 22429
rect 16025 22420 16037 22423
rect 15252 22392 16037 22420
rect 15252 22380 15258 22392
rect 16025 22389 16037 22392
rect 16071 22389 16083 22423
rect 18598 22420 18604 22432
rect 18559 22392 18604 22420
rect 16025 22383 16083 22389
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 19444 22429 19472 22732
rect 21082 22720 21088 22732
rect 21140 22760 21146 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 21140 22732 21189 22760
rect 21140 22720 21146 22732
rect 21177 22729 21189 22732
rect 21223 22729 21235 22763
rect 21177 22723 21235 22729
rect 21266 22720 21272 22772
rect 21324 22760 21330 22772
rect 22573 22763 22631 22769
rect 22573 22760 22585 22763
rect 21324 22732 22585 22760
rect 21324 22720 21330 22732
rect 22573 22729 22585 22732
rect 22619 22729 22631 22763
rect 22573 22723 22631 22729
rect 22741 22763 22799 22769
rect 22741 22729 22753 22763
rect 22787 22729 22799 22763
rect 22741 22723 22799 22729
rect 25041 22763 25099 22769
rect 25041 22729 25053 22763
rect 25087 22760 25099 22763
rect 27338 22760 27344 22772
rect 25087 22732 27344 22760
rect 25087 22729 25099 22732
rect 25041 22723 25099 22729
rect 20622 22692 20628 22704
rect 19536 22664 20628 22692
rect 19536 22633 19564 22664
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22593 19579 22627
rect 19521 22587 19579 22593
rect 20070 22584 20076 22636
rect 20128 22624 20134 22636
rect 20456 22633 20484 22664
rect 20622 22652 20628 22664
rect 20680 22692 20686 22704
rect 22094 22692 22100 22704
rect 20680 22664 22100 22692
rect 20680 22652 20686 22664
rect 22094 22652 22100 22664
rect 22152 22692 22158 22704
rect 22152 22664 22324 22692
rect 22152 22652 22158 22664
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 20128 22596 20177 22624
rect 20128 22584 20134 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22593 20499 22627
rect 20898 22624 20904 22636
rect 20441 22587 20499 22593
rect 20548 22596 20904 22624
rect 20349 22559 20407 22565
rect 20349 22525 20361 22559
rect 20395 22556 20407 22559
rect 20548 22556 20576 22596
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 21048 22596 21097 22624
rect 21048 22584 21054 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 21085 22587 21143 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 21818 22584 21824 22636
rect 21876 22624 21882 22636
rect 22296 22624 22324 22664
rect 22370 22652 22376 22704
rect 22428 22692 22434 22704
rect 22756 22692 22784 22723
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 28810 22760 28816 22772
rect 28771 22732 28816 22760
rect 28810 22720 28816 22732
rect 28868 22720 28874 22772
rect 29730 22760 29736 22772
rect 29691 22732 29736 22760
rect 29730 22720 29736 22732
rect 29788 22720 29794 22772
rect 29822 22720 29828 22772
rect 29880 22760 29886 22772
rect 30558 22760 30564 22772
rect 29880 22732 30564 22760
rect 29880 22720 29886 22732
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 30653 22763 30711 22769
rect 30653 22729 30665 22763
rect 30699 22760 30711 22763
rect 30742 22760 30748 22772
rect 30699 22732 30748 22760
rect 30699 22729 30711 22732
rect 30653 22723 30711 22729
rect 30742 22720 30748 22732
rect 30800 22720 30806 22772
rect 32217 22763 32275 22769
rect 32217 22729 32229 22763
rect 32263 22760 32275 22763
rect 32398 22760 32404 22772
rect 32263 22732 32404 22760
rect 32263 22729 32275 22732
rect 32217 22723 32275 22729
rect 32398 22720 32404 22732
rect 32456 22720 32462 22772
rect 25866 22692 25872 22704
rect 22428 22664 22473 22692
rect 22572 22664 22784 22692
rect 23308 22664 24164 22692
rect 22428 22652 22434 22664
rect 22572 22624 22600 22664
rect 23308 22633 23336 22664
rect 21876 22596 22232 22624
rect 22296 22596 22600 22624
rect 23293 22627 23351 22633
rect 21876 22584 21882 22596
rect 20395 22528 20576 22556
rect 21284 22556 21312 22584
rect 22204 22556 22232 22596
rect 23293 22593 23305 22627
rect 23339 22593 23351 22627
rect 23293 22587 23351 22593
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 23308 22556 23336 22587
rect 21284 22528 22094 22556
rect 22204 22528 23336 22556
rect 20395 22525 20407 22528
rect 20349 22519 20407 22525
rect 19705 22491 19763 22497
rect 19705 22457 19717 22491
rect 19751 22488 19763 22491
rect 20254 22488 20260 22500
rect 19751 22460 20260 22488
rect 19751 22457 19763 22460
rect 19705 22451 19763 22457
rect 20254 22448 20260 22460
rect 20312 22448 20318 22500
rect 20625 22491 20683 22497
rect 20625 22488 20637 22491
rect 20364 22460 20637 22488
rect 19429 22423 19487 22429
rect 19429 22389 19441 22423
rect 19475 22389 19487 22423
rect 19429 22383 19487 22389
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 20364 22420 20392 22460
rect 20625 22457 20637 22460
rect 20671 22457 20683 22491
rect 22066 22488 22094 22528
rect 23842 22488 23848 22500
rect 22066 22460 23848 22488
rect 20625 22451 20683 22457
rect 23842 22448 23848 22460
rect 23900 22448 23906 22500
rect 24044 22488 24072 22587
rect 24136 22556 24164 22664
rect 24228 22664 25872 22692
rect 24228 22633 24256 22664
rect 25866 22652 25872 22664
rect 25924 22652 25930 22704
rect 27522 22692 27528 22704
rect 27483 22664 27528 22692
rect 27522 22652 27528 22664
rect 27580 22692 27586 22704
rect 30098 22692 30104 22704
rect 27580 22664 28764 22692
rect 30059 22664 30104 22692
rect 27580 22652 27586 22664
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24946 22624 24952 22636
rect 24907 22596 24952 22624
rect 24213 22587 24271 22593
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 25593 22627 25651 22633
rect 25593 22593 25605 22627
rect 25639 22624 25651 22627
rect 26142 22624 26148 22636
rect 25639 22596 26148 22624
rect 25639 22593 25651 22596
rect 25593 22587 25651 22593
rect 26142 22584 26148 22596
rect 26200 22584 26206 22636
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22624 27767 22627
rect 27798 22624 27804 22636
rect 27755 22596 27804 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 27798 22584 27804 22596
rect 27856 22584 27862 22636
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 25498 22556 25504 22568
rect 24136 22528 25504 22556
rect 25498 22516 25504 22528
rect 25556 22556 25562 22568
rect 25869 22559 25927 22565
rect 25869 22556 25881 22559
rect 25556 22528 25881 22556
rect 25556 22516 25562 22528
rect 25869 22525 25881 22528
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 26050 22516 26056 22568
rect 26108 22556 26114 22568
rect 28000 22556 28028 22587
rect 28074 22584 28080 22636
rect 28132 22624 28138 22636
rect 28442 22624 28448 22636
rect 28132 22596 28448 22624
rect 28132 22584 28138 22596
rect 28442 22584 28448 22596
rect 28500 22624 28506 22636
rect 28736 22633 28764 22664
rect 30098 22652 30104 22664
rect 30156 22652 30162 22704
rect 32030 22652 32036 22704
rect 32088 22692 32094 22704
rect 32585 22695 32643 22701
rect 32585 22692 32597 22695
rect 32088 22664 32597 22692
rect 32088 22652 32094 22664
rect 32585 22661 32597 22664
rect 32631 22692 32643 22695
rect 32766 22692 32772 22704
rect 32631 22664 32772 22692
rect 32631 22661 32643 22664
rect 32585 22655 32643 22661
rect 32766 22652 32772 22664
rect 32824 22652 32830 22704
rect 32858 22652 32864 22704
rect 32916 22692 32922 22704
rect 33566 22695 33624 22701
rect 33566 22692 33578 22695
rect 32916 22664 33578 22692
rect 32916 22652 32922 22664
rect 33566 22661 33578 22664
rect 33612 22661 33624 22695
rect 33566 22655 33624 22661
rect 28537 22627 28595 22633
rect 28537 22624 28549 22627
rect 28500 22596 28549 22624
rect 28500 22584 28506 22596
rect 28537 22593 28549 22596
rect 28583 22593 28595 22627
rect 28537 22587 28595 22593
rect 28721 22627 28779 22633
rect 28721 22593 28733 22627
rect 28767 22593 28779 22627
rect 29914 22624 29920 22636
rect 29875 22596 29920 22624
rect 28721 22587 28779 22593
rect 29914 22584 29920 22596
rect 29972 22584 29978 22636
rect 30193 22627 30251 22633
rect 30193 22593 30205 22627
rect 30239 22624 30251 22627
rect 30239 22596 30328 22624
rect 30239 22593 30251 22596
rect 30193 22587 30251 22593
rect 30300 22568 30328 22596
rect 30834 22584 30840 22636
rect 30892 22633 30898 22636
rect 30892 22627 30941 22633
rect 30892 22593 30895 22627
rect 30929 22593 30941 22627
rect 31015 22624 31021 22636
rect 30976 22596 31021 22624
rect 30892 22587 30941 22593
rect 30892 22584 30898 22587
rect 31015 22584 31021 22596
rect 31073 22584 31079 22636
rect 31110 22584 31116 22636
rect 31168 22624 31174 22636
rect 31297 22627 31355 22633
rect 31168 22596 31213 22624
rect 31168 22584 31174 22596
rect 31297 22593 31309 22627
rect 31343 22593 31355 22627
rect 31297 22587 31355 22593
rect 26108 22528 28028 22556
rect 26108 22516 26114 22528
rect 30282 22516 30288 22568
rect 30340 22516 30346 22568
rect 30742 22516 30748 22568
rect 30800 22556 30806 22568
rect 31312 22556 31340 22587
rect 31754 22584 31760 22636
rect 31812 22624 31818 22636
rect 32306 22624 32312 22636
rect 31812 22596 32312 22624
rect 31812 22584 31818 22596
rect 32306 22584 32312 22596
rect 32364 22624 32370 22636
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 32364 22596 32413 22624
rect 32364 22584 32370 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32674 22624 32680 22636
rect 32635 22596 32680 22624
rect 32401 22587 32459 22593
rect 32674 22584 32680 22596
rect 32732 22584 32738 22636
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33321 22627 33379 22633
rect 33321 22624 33333 22627
rect 33192 22596 33333 22624
rect 33192 22584 33198 22596
rect 33321 22593 33333 22596
rect 33367 22624 33379 22627
rect 33410 22624 33416 22636
rect 33367 22596 33416 22624
rect 33367 22593 33379 22596
rect 33321 22587 33379 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 33226 22556 33232 22568
rect 30800 22528 33232 22556
rect 30800 22516 30806 22528
rect 33226 22516 33232 22528
rect 33284 22516 33290 22568
rect 25682 22488 25688 22500
rect 24044 22460 25688 22488
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 27798 22488 27804 22500
rect 27759 22460 27804 22488
rect 27798 22448 27804 22460
rect 27856 22448 27862 22500
rect 27890 22448 27896 22500
rect 27948 22488 27954 22500
rect 27948 22460 27993 22488
rect 27948 22448 27954 22460
rect 19576 22392 20392 22420
rect 20441 22423 20499 22429
rect 19576 22380 19582 22392
rect 20441 22389 20453 22423
rect 20487 22420 20499 22423
rect 20714 22420 20720 22432
rect 20487 22392 20720 22420
rect 20487 22389 20499 22392
rect 20441 22383 20499 22389
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 22554 22420 22560 22432
rect 22515 22392 22560 22420
rect 22554 22380 22560 22392
rect 22612 22380 22618 22432
rect 23385 22423 23443 22429
rect 23385 22389 23397 22423
rect 23431 22420 23443 22423
rect 23750 22420 23756 22432
rect 23431 22392 23756 22420
rect 23431 22389 23443 22392
rect 23385 22383 23443 22389
rect 23750 22380 23756 22392
rect 23808 22380 23814 22432
rect 24121 22423 24179 22429
rect 24121 22389 24133 22423
rect 24167 22420 24179 22423
rect 25958 22420 25964 22432
rect 24167 22392 25964 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 25958 22380 25964 22392
rect 26016 22380 26022 22432
rect 33318 22380 33324 22432
rect 33376 22420 33382 22432
rect 34701 22423 34759 22429
rect 34701 22420 34713 22423
rect 33376 22392 34713 22420
rect 33376 22380 33382 22392
rect 34701 22389 34713 22392
rect 34747 22389 34759 22423
rect 34701 22383 34759 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 17126 22176 17132 22228
rect 17184 22216 17190 22228
rect 17589 22219 17647 22225
rect 17589 22216 17601 22219
rect 17184 22188 17601 22216
rect 17184 22176 17190 22188
rect 17589 22185 17601 22188
rect 17635 22185 17647 22219
rect 19518 22216 19524 22228
rect 17589 22179 17647 22185
rect 17696 22188 19524 22216
rect 12434 22148 12440 22160
rect 12176 22120 12440 22148
rect 12176 22012 12204 22120
rect 12434 22108 12440 22120
rect 12492 22108 12498 22160
rect 13541 22151 13599 22157
rect 13541 22148 13553 22151
rect 13096 22120 13553 22148
rect 13096 22080 13124 22120
rect 13541 22117 13553 22120
rect 13587 22117 13599 22151
rect 17696 22148 17724 22188
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 19889 22219 19947 22225
rect 19889 22185 19901 22219
rect 19935 22216 19947 22219
rect 19978 22216 19984 22228
rect 19935 22188 19984 22216
rect 19935 22185 19947 22188
rect 19889 22179 19947 22185
rect 19978 22176 19984 22188
rect 20036 22216 20042 22228
rect 21266 22216 21272 22228
rect 20036 22188 21272 22216
rect 20036 22176 20042 22188
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 25590 22216 25596 22228
rect 24452 22188 25596 22216
rect 24452 22176 24458 22188
rect 25590 22176 25596 22188
rect 25648 22176 25654 22228
rect 25685 22219 25743 22225
rect 25685 22185 25697 22219
rect 25731 22216 25743 22219
rect 25958 22216 25964 22228
rect 25731 22188 25964 22216
rect 25731 22185 25743 22188
rect 25685 22179 25743 22185
rect 25958 22176 25964 22188
rect 26016 22176 26022 22228
rect 27798 22216 27804 22228
rect 27759 22188 27804 22216
rect 27798 22176 27804 22188
rect 27856 22216 27862 22228
rect 28442 22216 28448 22228
rect 27856 22188 28448 22216
rect 27856 22176 27862 22188
rect 28442 22176 28448 22188
rect 28500 22216 28506 22228
rect 28813 22219 28871 22225
rect 28813 22216 28825 22219
rect 28500 22188 28825 22216
rect 28500 22176 28506 22188
rect 28813 22185 28825 22188
rect 28859 22185 28871 22219
rect 29638 22216 29644 22228
rect 29599 22188 29644 22216
rect 28813 22179 28871 22185
rect 29638 22176 29644 22188
rect 29696 22176 29702 22228
rect 30285 22219 30343 22225
rect 30285 22185 30297 22219
rect 30331 22216 30343 22219
rect 30374 22216 30380 22228
rect 30331 22188 30380 22216
rect 30331 22185 30343 22188
rect 30285 22179 30343 22185
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 33318 22176 33324 22228
rect 33376 22216 33382 22228
rect 33597 22219 33655 22225
rect 33597 22216 33609 22219
rect 33376 22188 33609 22216
rect 33376 22176 33382 22188
rect 33597 22185 33609 22188
rect 33643 22185 33655 22219
rect 33597 22179 33655 22185
rect 13541 22111 13599 22117
rect 16408 22120 17724 22148
rect 14458 22080 14464 22092
rect 12360 22052 13124 22080
rect 13188 22052 14464 22080
rect 12360 22021 12388 22052
rect 12253 22015 12311 22021
rect 12253 22012 12265 22015
rect 12176 21984 12265 22012
rect 12253 21981 12265 21984
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 12989 22015 13047 22021
rect 12989 21981 13001 22015
rect 13035 22012 13047 22015
rect 13078 22012 13084 22024
rect 13035 21984 13084 22012
rect 13035 21981 13047 21984
rect 12989 21975 13047 21981
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13188 22021 13216 22052
rect 14458 22040 14464 22052
rect 14516 22040 14522 22092
rect 15028 22066 15424 22094
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 21981 13231 22015
rect 13354 22012 13360 22024
rect 13315 21984 13360 22012
rect 13173 21975 13231 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 14829 22015 14887 22021
rect 14829 21981 14841 22015
rect 14875 22012 14887 22015
rect 15028 22012 15056 22066
rect 14875 21984 15056 22012
rect 15197 22015 15255 22021
rect 14875 21981 14887 21984
rect 14829 21975 14887 21981
rect 15197 21981 15209 22015
rect 15243 22012 15255 22015
rect 15286 22012 15292 22024
rect 15243 21984 15292 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 15396 22012 15424 22066
rect 16408 22080 16436 22120
rect 19334 22108 19340 22160
rect 19392 22148 19398 22160
rect 20162 22148 20168 22160
rect 19392 22120 20168 22148
rect 19392 22108 19398 22120
rect 20162 22108 20168 22120
rect 20220 22108 20226 22160
rect 26970 22148 26976 22160
rect 25306 22120 26976 22148
rect 16485 22083 16543 22089
rect 16485 22080 16497 22083
rect 16408 22052 16497 22080
rect 16485 22049 16497 22052
rect 16531 22049 16543 22083
rect 16485 22043 16543 22049
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 16816 22052 17264 22080
rect 16816 22040 16822 22052
rect 15562 22012 15568 22024
rect 15396 21984 15568 22012
rect 15562 21972 15568 21984
rect 15620 22012 15626 22024
rect 16206 22012 16212 22024
rect 15620 21984 15976 22012
rect 16167 21984 16212 22012
rect 15620 21972 15626 21984
rect 13265 21947 13323 21953
rect 13265 21913 13277 21947
rect 13311 21944 13323 21947
rect 14274 21944 14280 21956
rect 13311 21916 14280 21944
rect 13311 21913 13323 21916
rect 13265 21907 13323 21913
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 15013 21947 15071 21953
rect 15013 21913 15025 21947
rect 15059 21913 15071 21947
rect 15013 21907 15071 21913
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 13446 21876 13452 21888
rect 12575 21848 13452 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 15028 21876 15056 21907
rect 15102 21904 15108 21956
rect 15160 21944 15166 21956
rect 15948 21944 15976 21984
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 17236 22021 17264 22052
rect 18138 22040 18144 22092
rect 18196 22080 18202 22092
rect 18417 22083 18475 22089
rect 18417 22080 18429 22083
rect 18196 22052 18429 22080
rect 18196 22040 18202 22052
rect 18417 22049 18429 22052
rect 18463 22049 18475 22083
rect 20898 22080 20904 22092
rect 20859 22052 20904 22080
rect 18417 22043 18475 22049
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 24578 22040 24584 22092
rect 24636 22080 24642 22092
rect 25306 22089 25334 22120
rect 26970 22108 26976 22120
rect 27028 22148 27034 22160
rect 29546 22148 29552 22160
rect 27028 22120 29552 22148
rect 27028 22108 27034 22120
rect 29546 22108 29552 22120
rect 29604 22108 29610 22160
rect 29656 22148 29684 22176
rect 29656 22120 30604 22148
rect 25133 22083 25191 22089
rect 25133 22080 25145 22083
rect 24636 22052 25145 22080
rect 24636 22040 24642 22052
rect 25133 22049 25145 22052
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 25291 22083 25349 22089
rect 25291 22049 25303 22083
rect 25337 22049 25349 22083
rect 25498 22080 25504 22092
rect 25459 22052 25504 22080
rect 25291 22043 25349 22049
rect 17037 22015 17095 22021
rect 17037 22012 17049 22015
rect 16408 21984 17049 22012
rect 16408 21944 16436 21984
rect 17037 21981 17049 21984
rect 17083 21981 17095 22015
rect 17037 21975 17095 21981
rect 17221 22015 17279 22021
rect 17221 21981 17233 22015
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 17310 21944 17316 21956
rect 15160 21916 15205 21944
rect 15304 21916 15884 21944
rect 15948 21916 16436 21944
rect 17271 21916 17316 21944
rect 15160 21904 15166 21916
rect 15304 21876 15332 21916
rect 15028 21848 15332 21876
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 15856 21885 15884 21916
rect 17310 21904 17316 21916
rect 17368 21904 17374 21956
rect 15841 21879 15899 21885
rect 15436 21848 15481 21876
rect 15436 21836 15442 21848
rect 15841 21845 15853 21879
rect 15887 21845 15899 21879
rect 16298 21876 16304 21888
rect 16259 21848 16304 21876
rect 15841 21839 15899 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 16482 21836 16488 21888
rect 16540 21876 16546 21888
rect 17420 21876 17448 21975
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18325 22015 18383 22021
rect 18325 22012 18337 22015
rect 18288 21984 18337 22012
rect 18288 21972 18294 21984
rect 18325 21981 18337 21984
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 19334 22012 19340 22024
rect 18555 21984 19340 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 20165 22015 20223 22021
rect 20165 21981 20177 22015
rect 20211 22012 20223 22015
rect 20530 22012 20536 22024
rect 20211 21984 20536 22012
rect 20211 21981 20223 21984
rect 20165 21975 20223 21981
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 22097 22015 22155 22021
rect 20680 21984 20725 22012
rect 20680 21972 20686 21984
rect 22097 21981 22109 22015
rect 22143 22012 22155 22015
rect 23106 22012 23112 22024
rect 22143 21984 23112 22012
rect 22143 21981 22155 21984
rect 22097 21975 22155 21981
rect 23106 21972 23112 21984
rect 23164 22012 23170 22024
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 23164 21984 24685 22012
rect 23164 21972 23170 21984
rect 24673 21981 24685 21984
rect 24719 22012 24731 22015
rect 24854 22012 24860 22024
rect 24719 21984 24860 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 19705 21947 19763 21953
rect 19705 21913 19717 21947
rect 19751 21944 19763 21947
rect 22364 21947 22422 21953
rect 19751 21916 22094 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 16540 21848 17448 21876
rect 19889 21879 19947 21885
rect 16540 21836 16546 21848
rect 19889 21845 19901 21879
rect 19935 21876 19947 21879
rect 19978 21876 19984 21888
rect 19935 21848 19984 21876
rect 19935 21845 19947 21848
rect 19889 21839 19947 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 22066 21876 22094 21916
rect 22364 21913 22376 21947
rect 22410 21944 22422 21947
rect 23014 21944 23020 21956
rect 22410 21916 23020 21944
rect 22410 21913 22422 21916
rect 22364 21907 22422 21913
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 24210 21944 24216 21956
rect 23124 21916 24216 21944
rect 23124 21876 23152 21916
rect 24210 21904 24216 21916
rect 24268 21904 24274 21956
rect 24486 21944 24492 21956
rect 24447 21916 24492 21944
rect 24486 21904 24492 21916
rect 24544 21904 24550 21956
rect 23474 21876 23480 21888
rect 22066 21848 23152 21876
rect 23435 21848 23480 21876
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 25148 21876 25176 22043
rect 25498 22040 25504 22052
rect 25556 22040 25562 22092
rect 28166 22040 28172 22092
rect 28224 22080 28230 22092
rect 29825 22083 29883 22089
rect 28224 22052 28672 22080
rect 28224 22040 28230 22052
rect 25866 21972 25872 22024
rect 25924 22012 25930 22024
rect 25924 21984 26188 22012
rect 25924 21972 25930 21984
rect 26160 21953 26188 21984
rect 26234 21972 26240 22024
rect 26292 22012 26298 22024
rect 26421 22015 26479 22021
rect 26421 22012 26433 22015
rect 26292 21984 26433 22012
rect 26292 21972 26298 21984
rect 26421 21981 26433 21984
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 26697 22015 26755 22021
rect 26697 21981 26709 22015
rect 26743 22012 26755 22015
rect 27341 22015 27399 22021
rect 27341 22012 27353 22015
rect 26743 21984 27353 22012
rect 26743 21981 26755 21984
rect 26697 21975 26755 21981
rect 27341 21981 27353 21984
rect 27387 21981 27399 22015
rect 27706 22012 27712 22024
rect 27667 21984 27712 22012
rect 27341 21975 27399 21981
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 27890 21972 27896 22024
rect 27948 22012 27954 22024
rect 27985 22015 28043 22021
rect 27985 22012 27997 22015
rect 27948 21984 27997 22012
rect 27948 21972 27954 21984
rect 27985 21981 27997 21984
rect 28031 22012 28043 22015
rect 28031 21984 28304 22012
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 26145 21947 26203 21953
rect 26145 21913 26157 21947
rect 26191 21913 26203 21947
rect 26145 21907 26203 21913
rect 26326 21876 26332 21888
rect 25148 21848 26332 21876
rect 26326 21836 26332 21848
rect 26384 21836 26390 21888
rect 26510 21876 26516 21888
rect 26471 21848 26516 21876
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 27522 21876 27528 21888
rect 27483 21848 27528 21876
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 28276 21876 28304 21984
rect 28350 21972 28356 22024
rect 28408 22012 28414 22024
rect 28445 22015 28503 22021
rect 28445 22012 28457 22015
rect 28408 21984 28457 22012
rect 28408 21972 28414 21984
rect 28445 21981 28457 21984
rect 28491 21981 28503 22015
rect 28445 21975 28503 21981
rect 28644 21953 28672 22052
rect 29825 22049 29837 22083
rect 29871 22080 29883 22083
rect 29914 22080 29920 22092
rect 29871 22052 29920 22080
rect 29871 22049 29883 22052
rect 29825 22043 29883 22049
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 30190 22040 30196 22092
rect 30248 22080 30254 22092
rect 30248 22052 30512 22080
rect 30248 22040 30254 22052
rect 29549 22015 29607 22021
rect 29549 21981 29561 22015
rect 29595 22012 29607 22015
rect 29638 22012 29644 22024
rect 29595 21984 29644 22012
rect 29595 21981 29607 21984
rect 29549 21975 29607 21981
rect 29638 21972 29644 21984
rect 29696 21972 29702 22024
rect 30282 22012 30288 22024
rect 30243 21984 30288 22012
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 30484 22021 30512 22052
rect 30469 22015 30527 22021
rect 30469 21981 30481 22015
rect 30515 21981 30527 22015
rect 30576 22012 30604 22120
rect 32490 22108 32496 22160
rect 32548 22148 32554 22160
rect 32548 22120 32812 22148
rect 32548 22108 32554 22120
rect 31205 22083 31263 22089
rect 31205 22049 31217 22083
rect 31251 22080 31263 22083
rect 32508 22080 32536 22108
rect 32674 22080 32680 22092
rect 31251 22052 32536 22080
rect 32635 22052 32680 22080
rect 31251 22049 31263 22052
rect 31205 22043 31263 22049
rect 32674 22040 32680 22052
rect 32732 22040 32738 22092
rect 32784 22089 32812 22120
rect 32769 22083 32827 22089
rect 32769 22049 32781 22083
rect 32815 22080 32827 22083
rect 33318 22080 33324 22092
rect 32815 22052 33324 22080
rect 32815 22049 32827 22052
rect 32769 22043 32827 22049
rect 33318 22040 33324 22052
rect 33376 22040 33382 22092
rect 33781 22083 33839 22089
rect 33781 22049 33793 22083
rect 33827 22080 33839 22083
rect 34790 22080 34796 22092
rect 33827 22052 34796 22080
rect 33827 22049 33839 22052
rect 33781 22043 33839 22049
rect 34790 22040 34796 22052
rect 34848 22040 34854 22092
rect 30929 22015 30987 22021
rect 30929 22012 30941 22015
rect 30576 21984 30941 22012
rect 30469 21975 30527 21981
rect 30929 21981 30941 21984
rect 30975 22012 30987 22015
rect 31294 22012 31300 22024
rect 30975 21984 31300 22012
rect 30975 21981 30987 21984
rect 30929 21975 30987 21981
rect 31294 21972 31300 21984
rect 31352 21972 31358 22024
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 32401 22015 32459 22021
rect 32401 22012 32413 22015
rect 32180 21984 32413 22012
rect 32180 21972 32186 21984
rect 32401 21981 32413 21984
rect 32447 21981 32459 22015
rect 32401 21975 32459 21981
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 32585 22015 32643 22021
rect 32585 22012 32597 22015
rect 32548 21984 32597 22012
rect 32548 21972 32554 21984
rect 32585 21981 32597 21984
rect 32631 21981 32643 22015
rect 32585 21975 32643 21981
rect 32953 22015 33011 22021
rect 32953 21981 32965 22015
rect 32999 22012 33011 22015
rect 33042 22012 33048 22024
rect 32999 21984 33048 22012
rect 32999 21981 33011 21984
rect 32953 21975 33011 21981
rect 33042 21972 33048 21984
rect 33100 22012 33106 22024
rect 33873 22015 33931 22021
rect 33100 21984 33640 22012
rect 33100 21972 33106 21984
rect 33612 21956 33640 21984
rect 33873 21981 33885 22015
rect 33919 22012 33931 22015
rect 34698 22012 34704 22024
rect 33919 21984 34704 22012
rect 33919 21981 33931 21984
rect 33873 21975 33931 21981
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 28629 21947 28687 21953
rect 28629 21913 28641 21947
rect 28675 21913 28687 21947
rect 29822 21944 29828 21956
rect 29783 21916 29828 21944
rect 28629 21907 28687 21913
rect 29822 21904 29828 21916
rect 29880 21904 29886 21956
rect 33594 21944 33600 21956
rect 31496 21916 33272 21944
rect 33555 21916 33600 21944
rect 31496 21876 31524 21916
rect 33134 21876 33140 21888
rect 28276 21848 31524 21876
rect 33095 21848 33140 21876
rect 33134 21836 33140 21848
rect 33192 21836 33198 21888
rect 33244 21876 33272 21916
rect 33594 21904 33600 21916
rect 33652 21904 33658 21956
rect 34057 21879 34115 21885
rect 34057 21876 34069 21879
rect 33244 21848 34069 21876
rect 34057 21845 34069 21848
rect 34103 21845 34115 21879
rect 34057 21839 34115 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 16482 21672 16488 21684
rect 15344 21644 16488 21672
rect 15344 21632 15350 21644
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 17129 21675 17187 21681
rect 17129 21641 17141 21675
rect 17175 21672 17187 21675
rect 17770 21672 17776 21684
rect 17175 21644 17776 21672
rect 17175 21641 17187 21644
rect 17129 21635 17187 21641
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20622 21672 20628 21684
rect 20220 21644 20628 21672
rect 20220 21632 20226 21644
rect 20622 21632 20628 21644
rect 20680 21672 20686 21684
rect 22189 21675 22247 21681
rect 22189 21672 22201 21675
rect 20680 21644 22201 21672
rect 20680 21632 20686 21644
rect 22189 21641 22201 21644
rect 22235 21641 22247 21675
rect 22189 21635 22247 21641
rect 22925 21675 22983 21681
rect 22925 21641 22937 21675
rect 22971 21672 22983 21675
rect 24302 21672 24308 21684
rect 22971 21644 24308 21672
rect 22971 21641 22983 21644
rect 22925 21635 22983 21641
rect 24302 21632 24308 21644
rect 24360 21632 24366 21684
rect 24673 21675 24731 21681
rect 24673 21641 24685 21675
rect 24719 21672 24731 21675
rect 25406 21672 25412 21684
rect 24719 21644 25412 21672
rect 24719 21641 24731 21644
rect 24673 21635 24731 21641
rect 25406 21632 25412 21644
rect 25464 21672 25470 21684
rect 26050 21672 26056 21684
rect 25464 21644 26056 21672
rect 25464 21632 25470 21644
rect 26050 21632 26056 21644
rect 26108 21632 26114 21684
rect 26970 21632 26976 21684
rect 27028 21672 27034 21684
rect 31202 21672 31208 21684
rect 27028 21644 28304 21672
rect 31163 21644 31208 21672
rect 27028 21632 27034 21644
rect 15102 21564 15108 21616
rect 15160 21604 15166 21616
rect 16298 21604 16304 21616
rect 15160 21576 16304 21604
rect 15160 21564 15166 21576
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 21818 21604 21824 21616
rect 21779 21576 21824 21604
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 22002 21564 22008 21616
rect 22060 21613 22066 21616
rect 22060 21607 22079 21613
rect 22067 21573 22079 21607
rect 22060 21567 22079 21573
rect 22060 21564 22066 21567
rect 23014 21564 23020 21616
rect 23072 21604 23078 21616
rect 23293 21607 23351 21613
rect 23293 21604 23305 21607
rect 23072 21576 23305 21604
rect 23072 21564 23078 21576
rect 23293 21573 23305 21576
rect 23339 21573 23351 21607
rect 25590 21604 25596 21616
rect 23293 21567 23351 21573
rect 23400 21576 25596 21604
rect 12802 21536 12808 21548
rect 12763 21508 12808 21536
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 13078 21545 13084 21548
rect 13072 21499 13084 21545
rect 13136 21536 13142 21548
rect 13136 21508 13172 21536
rect 13078 21496 13084 21499
rect 13136 21496 13142 21508
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 14993 21539 15051 21545
rect 14993 21536 15005 21539
rect 14884 21508 15005 21536
rect 14884 21496 14890 21508
rect 14993 21505 15005 21508
rect 15039 21505 15051 21539
rect 14993 21499 15051 21505
rect 15746 21496 15752 21548
rect 15804 21536 15810 21548
rect 16761 21539 16819 21545
rect 16761 21536 16773 21539
rect 15804 21508 16773 21536
rect 15804 21496 15810 21508
rect 16761 21505 16773 21508
rect 16807 21505 16819 21539
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 16761 21499 16819 21505
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18305 21539 18363 21545
rect 18305 21536 18317 21539
rect 18196 21508 18317 21536
rect 18196 21496 18202 21508
rect 18305 21505 18317 21508
rect 18351 21505 18363 21539
rect 20438 21536 20444 21548
rect 20399 21508 20444 21536
rect 18305 21499 18363 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 20714 21536 20720 21548
rect 20675 21508 20720 21536
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 22554 21536 22560 21548
rect 22020 21508 22560 21536
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 13872 21440 14749 21468
rect 13872 21428 13878 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 14185 21335 14243 21341
rect 14185 21301 14197 21335
rect 14231 21332 14243 21335
rect 14274 21332 14280 21344
rect 14231 21304 14280 21332
rect 14231 21301 14243 21304
rect 14185 21295 14243 21301
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14752 21332 14780 21431
rect 16390 21360 16396 21412
rect 16448 21400 16454 21412
rect 18064 21400 18092 21431
rect 16448 21372 18092 21400
rect 16448 21360 16454 21372
rect 15470 21332 15476 21344
rect 14752 21304 15476 21332
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16117 21335 16175 21341
rect 16117 21301 16129 21335
rect 16163 21332 16175 21335
rect 17310 21332 17316 21344
rect 16163 21304 17316 21332
rect 16163 21301 16175 21304
rect 16117 21295 16175 21301
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 19429 21335 19487 21341
rect 19429 21332 19441 21335
rect 19300 21304 19441 21332
rect 19300 21292 19306 21304
rect 19429 21301 19441 21304
rect 19475 21332 19487 21335
rect 20990 21332 20996 21344
rect 19475 21304 20996 21332
rect 19475 21301 19487 21304
rect 19429 21295 19487 21301
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 22020 21341 22048 21508
rect 22554 21496 22560 21508
rect 22612 21536 22618 21548
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 22612 21508 22845 21536
rect 22612 21496 22618 21508
rect 22833 21505 22845 21508
rect 22879 21536 22891 21539
rect 23400 21536 23428 21576
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 25958 21564 25964 21616
rect 26016 21604 26022 21616
rect 26145 21607 26203 21613
rect 26145 21604 26157 21607
rect 26016 21576 26157 21604
rect 26016 21564 26022 21576
rect 26145 21573 26157 21576
rect 26191 21573 26203 21607
rect 26145 21567 26203 21573
rect 27157 21607 27215 21613
rect 27157 21573 27169 21607
rect 27203 21604 27215 21607
rect 27982 21604 27988 21616
rect 27203 21576 27988 21604
rect 27203 21573 27215 21576
rect 27157 21567 27215 21573
rect 27982 21564 27988 21576
rect 28040 21564 28046 21616
rect 22879 21508 23428 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 23474 21496 23480 21548
rect 23532 21536 23538 21548
rect 23753 21539 23811 21545
rect 23753 21536 23765 21539
rect 23532 21508 23765 21536
rect 23532 21496 23538 21508
rect 23753 21505 23765 21508
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21536 24639 21539
rect 24854 21536 24860 21548
rect 24627 21508 24860 21536
rect 24627 21505 24639 21508
rect 24581 21499 24639 21505
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21536 25467 21539
rect 25682 21536 25688 21548
rect 25455 21508 25688 21536
rect 25455 21505 25467 21508
rect 25409 21499 25467 21505
rect 25682 21496 25688 21508
rect 25740 21536 25746 21548
rect 26510 21536 26516 21548
rect 25740 21508 26516 21536
rect 25740 21496 25746 21508
rect 26510 21496 26516 21508
rect 26568 21496 26574 21548
rect 27522 21496 27528 21548
rect 27580 21536 27586 21548
rect 28276 21545 28304 21644
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 32125 21675 32183 21681
rect 32125 21641 32137 21675
rect 32171 21672 32183 21675
rect 32674 21672 32680 21684
rect 32171 21644 32680 21672
rect 32171 21641 32183 21644
rect 32125 21635 32183 21641
rect 32674 21632 32680 21644
rect 32732 21632 32738 21684
rect 33594 21632 33600 21684
rect 33652 21672 33658 21684
rect 34885 21675 34943 21681
rect 34885 21672 34897 21675
rect 33652 21644 34897 21672
rect 33652 21632 33658 21644
rect 34885 21641 34897 21644
rect 34931 21641 34943 21675
rect 34885 21635 34943 21641
rect 30469 21607 30527 21613
rect 30469 21573 30481 21607
rect 30515 21604 30527 21607
rect 30929 21607 30987 21613
rect 30929 21604 30941 21607
rect 30515 21576 30941 21604
rect 30515 21573 30527 21576
rect 30469 21567 30527 21573
rect 30929 21573 30941 21576
rect 30975 21573 30987 21607
rect 30929 21567 30987 21573
rect 31113 21607 31171 21613
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 31159 21576 32444 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 32416 21548 32444 21576
rect 33134 21564 33140 21616
rect 33192 21604 33198 21616
rect 33750 21607 33808 21613
rect 33750 21604 33762 21607
rect 33192 21576 33762 21604
rect 33192 21564 33198 21576
rect 33750 21573 33762 21576
rect 33796 21573 33808 21607
rect 33750 21567 33808 21573
rect 33870 21564 33876 21616
rect 33928 21604 33934 21616
rect 35621 21607 35679 21613
rect 35621 21604 35633 21607
rect 33928 21576 35633 21604
rect 33928 21564 33934 21576
rect 35621 21573 35633 21576
rect 35667 21573 35679 21607
rect 35621 21567 35679 21573
rect 28077 21539 28135 21545
rect 28077 21536 28089 21539
rect 27580 21508 28089 21536
rect 27580 21496 27586 21508
rect 28077 21505 28089 21508
rect 28123 21505 28135 21539
rect 28077 21499 28135 21505
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 28261 21539 28319 21545
rect 28261 21505 28273 21539
rect 28307 21505 28319 21539
rect 28442 21536 28448 21548
rect 28403 21508 28448 21536
rect 28261 21499 28319 21505
rect 23198 21468 23204 21480
rect 23159 21440 23204 21468
rect 23198 21428 23204 21440
rect 23256 21428 23262 21480
rect 25225 21471 25283 21477
rect 25225 21437 25237 21471
rect 25271 21468 25283 21471
rect 25958 21468 25964 21480
rect 25271 21440 25964 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 25958 21428 25964 21440
rect 26016 21428 26022 21480
rect 27706 21428 27712 21480
rect 27764 21468 27770 21480
rect 28184 21468 28212 21499
rect 28442 21496 28448 21508
rect 28500 21496 28506 21548
rect 29178 21536 29184 21548
rect 29139 21508 29184 21536
rect 29178 21496 29184 21508
rect 29236 21496 29242 21548
rect 29273 21539 29331 21545
rect 29273 21505 29285 21539
rect 29319 21505 29331 21539
rect 29273 21499 29331 21505
rect 29365 21539 29423 21545
rect 29365 21505 29377 21539
rect 29411 21505 29423 21539
rect 29546 21536 29552 21548
rect 29507 21508 29552 21536
rect 29365 21499 29423 21505
rect 29288 21468 29316 21499
rect 27764 21440 29316 21468
rect 29380 21468 29408 21499
rect 29546 21496 29552 21508
rect 29604 21496 29610 21548
rect 30006 21496 30012 21548
rect 30064 21536 30070 21548
rect 30190 21536 30196 21548
rect 30064 21508 30196 21536
rect 30064 21496 30070 21508
rect 30190 21496 30196 21508
rect 30248 21496 30254 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 31294 21536 31300 21548
rect 31251 21508 31300 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 31294 21496 31300 21508
rect 31352 21536 31358 21548
rect 32306 21536 32312 21548
rect 31352 21508 31754 21536
rect 32267 21508 32312 21536
rect 31352 21496 31358 21508
rect 29638 21468 29644 21480
rect 29380 21440 29644 21468
rect 27764 21428 27770 21440
rect 29638 21428 29644 21440
rect 29696 21468 29702 21480
rect 30098 21468 30104 21480
rect 29696 21440 30104 21468
rect 29696 21428 29702 21440
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 30469 21471 30527 21477
rect 30469 21437 30481 21471
rect 30515 21468 30527 21471
rect 30558 21468 30564 21480
rect 30515 21440 30564 21468
rect 30515 21437 30527 21440
rect 30469 21431 30527 21437
rect 30558 21428 30564 21440
rect 30616 21428 30622 21480
rect 23109 21403 23167 21409
rect 23109 21369 23121 21403
rect 23155 21400 23167 21403
rect 23658 21400 23664 21412
rect 23155 21372 23664 21400
rect 23155 21369 23167 21372
rect 23109 21363 23167 21369
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 24762 21360 24768 21412
rect 24820 21400 24826 21412
rect 26329 21403 26387 21409
rect 26329 21400 26341 21403
rect 24820 21372 26341 21400
rect 24820 21360 24826 21372
rect 26329 21369 26341 21372
rect 26375 21369 26387 21403
rect 26329 21363 26387 21369
rect 27341 21403 27399 21409
rect 27341 21369 27353 21403
rect 27387 21400 27399 21403
rect 27387 21372 28212 21400
rect 27387 21369 27399 21372
rect 27341 21363 27399 21369
rect 22005 21335 22063 21341
rect 22005 21301 22017 21335
rect 22051 21301 22063 21335
rect 23750 21332 23756 21344
rect 23711 21304 23756 21332
rect 22005 21295 22063 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 25314 21292 25320 21344
rect 25372 21332 25378 21344
rect 26142 21332 26148 21344
rect 25372 21304 26148 21332
rect 25372 21292 25378 21304
rect 26142 21292 26148 21304
rect 26200 21292 26206 21344
rect 27798 21332 27804 21344
rect 27759 21304 27804 21332
rect 27798 21292 27804 21304
rect 27856 21292 27862 21344
rect 28184 21332 28212 21372
rect 28718 21332 28724 21344
rect 28184 21304 28724 21332
rect 28718 21292 28724 21304
rect 28776 21292 28782 21344
rect 28905 21335 28963 21341
rect 28905 21301 28917 21335
rect 28951 21332 28963 21335
rect 28994 21332 29000 21344
rect 28951 21304 29000 21332
rect 28951 21301 28963 21304
rect 28905 21295 28963 21301
rect 28994 21292 29000 21304
rect 29052 21292 29058 21344
rect 29914 21292 29920 21344
rect 29972 21332 29978 21344
rect 30282 21332 30288 21344
rect 29972 21304 30288 21332
rect 29972 21292 29978 21304
rect 30282 21292 30288 21304
rect 30340 21292 30346 21344
rect 31726 21332 31754 21508
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 32398 21496 32404 21548
rect 32456 21536 32462 21548
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 32456 21508 32505 21536
rect 32456 21496 32462 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 32585 21539 32643 21545
rect 32585 21505 32597 21539
rect 32631 21536 32643 21539
rect 32858 21536 32864 21548
rect 32631 21508 32864 21536
rect 32631 21505 32643 21508
rect 32585 21499 32643 21505
rect 32306 21360 32312 21412
rect 32364 21400 32370 21412
rect 32600 21400 32628 21499
rect 32858 21496 32864 21508
rect 32916 21496 32922 21548
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 35345 21539 35403 21545
rect 35345 21536 35357 21539
rect 34848 21508 35357 21536
rect 34848 21496 34854 21508
rect 35345 21505 35357 21508
rect 35391 21505 35403 21539
rect 35345 21499 35403 21505
rect 33502 21468 33508 21480
rect 33463 21440 33508 21468
rect 33502 21428 33508 21440
rect 33560 21428 33566 21480
rect 35618 21468 35624 21480
rect 35579 21440 35624 21468
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 32364 21372 32628 21400
rect 32364 21360 32370 21372
rect 35437 21335 35495 21341
rect 35437 21332 35449 21335
rect 31726 21304 35449 21332
rect 35437 21301 35449 21304
rect 35483 21301 35495 21335
rect 35437 21295 35495 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13265 21131 13323 21137
rect 13265 21128 13277 21131
rect 13136 21100 13277 21128
rect 13136 21088 13142 21100
rect 13265 21097 13277 21100
rect 13311 21097 13323 21131
rect 13265 21091 13323 21097
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 14826 21128 14832 21140
rect 14783 21100 14832 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 15470 21088 15476 21140
rect 15528 21128 15534 21140
rect 15565 21131 15623 21137
rect 15565 21128 15577 21131
rect 15528 21100 15577 21128
rect 15528 21088 15534 21100
rect 15565 21097 15577 21100
rect 15611 21128 15623 21131
rect 16390 21128 16396 21140
rect 15611 21100 16396 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 19116 21100 19257 21128
rect 19116 21088 19122 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 19352 21100 19555 21128
rect 16574 21020 16580 21072
rect 16632 21060 16638 21072
rect 16942 21060 16948 21072
rect 16632 21032 16948 21060
rect 16632 21020 16638 21032
rect 16942 21020 16948 21032
rect 17000 21060 17006 21072
rect 19352 21060 19380 21100
rect 17000 21032 19380 21060
rect 19527 21060 19555 21100
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 20036 21100 20085 21128
rect 20036 21088 20042 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 20073 21091 20131 21097
rect 21818 21088 21824 21140
rect 21876 21128 21882 21140
rect 23750 21128 23756 21140
rect 21876 21100 23756 21128
rect 21876 21088 21882 21100
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 24765 21131 24823 21137
rect 24765 21097 24777 21131
rect 24811 21128 24823 21131
rect 25130 21128 25136 21140
rect 24811 21100 25136 21128
rect 24811 21097 24823 21100
rect 24765 21091 24823 21097
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 25774 21088 25780 21140
rect 25832 21128 25838 21140
rect 25832 21100 26372 21128
rect 25832 21088 25838 21100
rect 22646 21060 22652 21072
rect 19527 21032 22094 21060
rect 22607 21032 22652 21060
rect 17000 21020 17006 21032
rect 15102 20952 15108 21004
rect 15160 20992 15166 21004
rect 15160 20964 17172 20992
rect 15160 20952 15166 20964
rect 13446 20924 13452 20936
rect 13407 20896 13452 20924
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 15194 20924 15200 20936
rect 14967 20896 15200 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20924 15531 20927
rect 15562 20924 15568 20936
rect 15519 20896 15568 20924
rect 15519 20893 15531 20896
rect 15473 20887 15531 20893
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 16574 20924 16580 20936
rect 16535 20896 16580 20924
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 16758 20924 16764 20936
rect 16719 20896 16764 20924
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20924 17003 20927
rect 17034 20924 17040 20936
rect 16991 20896 17040 20924
rect 16991 20893 17003 20896
rect 16945 20887 17003 20893
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 16868 20856 16896 20887
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 17144 20933 17172 20964
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 19392 20964 20637 20992
rect 19392 20952 19398 20964
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 22066 20992 22094 21032
rect 22646 21020 22652 21032
rect 22704 21020 22710 21072
rect 22738 21020 22744 21072
rect 22796 21060 22802 21072
rect 23198 21060 23204 21072
rect 22796 21032 23204 21060
rect 22796 21020 22802 21032
rect 23198 21020 23204 21032
rect 23256 21020 23262 21072
rect 23290 21020 23296 21072
rect 23348 21060 23354 21072
rect 23477 21063 23535 21069
rect 23477 21060 23489 21063
rect 23348 21032 23489 21060
rect 23348 21020 23354 21032
rect 23477 21029 23489 21032
rect 23523 21029 23535 21063
rect 26344 21060 26372 21100
rect 26418 21088 26424 21140
rect 26476 21128 26482 21140
rect 26789 21131 26847 21137
rect 26789 21128 26801 21131
rect 26476 21100 26801 21128
rect 26476 21088 26482 21100
rect 26789 21097 26801 21100
rect 26835 21128 26847 21131
rect 27246 21128 27252 21140
rect 26835 21100 27252 21128
rect 26835 21097 26847 21100
rect 26789 21091 26847 21097
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 28258 21088 28264 21140
rect 28316 21128 28322 21140
rect 28353 21131 28411 21137
rect 28353 21128 28365 21131
rect 28316 21100 28365 21128
rect 28316 21088 28322 21100
rect 28353 21097 28365 21100
rect 28399 21097 28411 21131
rect 28353 21091 28411 21097
rect 28902 21088 28908 21140
rect 28960 21128 28966 21140
rect 29178 21128 29184 21140
rect 28960 21100 29184 21128
rect 28960 21088 28966 21100
rect 29178 21088 29184 21100
rect 29236 21088 29242 21140
rect 29270 21088 29276 21140
rect 29328 21128 29334 21140
rect 29549 21131 29607 21137
rect 29549 21128 29561 21131
rect 29328 21100 29561 21128
rect 29328 21088 29334 21100
rect 29549 21097 29561 21100
rect 29595 21097 29607 21131
rect 29549 21091 29607 21097
rect 29914 21088 29920 21140
rect 29972 21128 29978 21140
rect 30653 21131 30711 21137
rect 30653 21128 30665 21131
rect 29972 21100 30665 21128
rect 29972 21088 29978 21100
rect 30653 21097 30665 21100
rect 30699 21097 30711 21131
rect 30653 21091 30711 21097
rect 31665 21131 31723 21137
rect 31665 21097 31677 21131
rect 31711 21128 31723 21131
rect 32306 21128 32312 21140
rect 31711 21100 32312 21128
rect 31711 21097 31723 21100
rect 31665 21091 31723 21097
rect 32306 21088 32312 21100
rect 32364 21088 32370 21140
rect 32490 21088 32496 21140
rect 32548 21128 32554 21140
rect 33965 21131 34023 21137
rect 33965 21128 33977 21131
rect 32548 21100 33977 21128
rect 32548 21088 32554 21100
rect 33965 21097 33977 21100
rect 34011 21097 34023 21131
rect 33965 21091 34023 21097
rect 27617 21063 27675 21069
rect 27617 21060 27629 21063
rect 26344 21032 27629 21060
rect 23477 21023 23535 21029
rect 27617 21029 27629 21032
rect 27663 21060 27675 21063
rect 27706 21060 27712 21072
rect 27663 21032 27712 21060
rect 27663 21029 27675 21032
rect 27617 21023 27675 21029
rect 27706 21020 27712 21032
rect 27764 21020 27770 21072
rect 28810 21020 28816 21072
rect 28868 21060 28874 21072
rect 30190 21060 30196 21072
rect 28868 21032 30196 21060
rect 28868 21020 28874 21032
rect 30190 21020 30196 21032
rect 30248 21060 30254 21072
rect 31021 21063 31079 21069
rect 30248 21032 30788 21060
rect 30248 21020 30254 21032
rect 24854 20992 24860 21004
rect 22066 20964 24860 20992
rect 20625 20955 20683 20961
rect 17129 20927 17187 20933
rect 17129 20893 17141 20927
rect 17175 20893 17187 20927
rect 17129 20887 17187 20893
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 17359 20896 18245 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18414 20924 18420 20936
rect 18375 20896 18420 20924
rect 18233 20887 18291 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 19058 20924 19064 20936
rect 18555 20896 19064 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20924 19487 20927
rect 20070 20924 20076 20936
rect 19475 20896 20076 20924
rect 19475 20893 19487 20896
rect 19429 20887 19487 20893
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 22480 20933 22508 20964
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 26970 20952 26976 21004
rect 27028 20992 27034 21004
rect 27801 20995 27859 21001
rect 27801 20992 27813 20995
rect 27028 20964 27813 20992
rect 27028 20952 27034 20964
rect 27801 20961 27813 20964
rect 27847 20961 27859 20995
rect 27801 20955 27859 20961
rect 27890 20952 27896 21004
rect 27948 20992 27954 21004
rect 28546 20992 28672 21000
rect 27948 20972 28871 20992
rect 27948 20964 28574 20972
rect 28644 20964 28871 20972
rect 27948 20952 27954 20964
rect 21729 20927 21787 20933
rect 21729 20924 21741 20927
rect 20180 20896 21741 20924
rect 16080 20828 16896 20856
rect 16080 20816 16086 20828
rect 17678 20816 17684 20868
rect 17736 20856 17742 20868
rect 20180 20856 20208 20896
rect 21729 20893 21741 20896
rect 21775 20893 21787 20927
rect 21729 20887 21787 20893
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20924 21971 20927
rect 22465 20927 22523 20933
rect 21959 20896 22094 20924
rect 21959 20893 21971 20896
rect 21913 20887 21971 20893
rect 17736 20828 20208 20856
rect 20441 20859 20499 20865
rect 17736 20816 17742 20828
rect 20441 20825 20453 20859
rect 20487 20856 20499 20859
rect 21450 20856 21456 20868
rect 20487 20828 21456 20856
rect 20487 20825 20499 20828
rect 20441 20819 20499 20825
rect 21450 20816 21456 20828
rect 21508 20816 21514 20868
rect 22066 20856 22094 20896
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 23293 20927 23351 20933
rect 22465 20887 22523 20893
rect 22664 20896 23244 20924
rect 22664 20856 22692 20896
rect 22066 20828 22692 20856
rect 18046 20788 18052 20800
rect 18007 20760 18052 20788
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 21821 20791 21879 20797
rect 20588 20760 20633 20788
rect 20588 20748 20594 20760
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22186 20788 22192 20800
rect 21867 20760 22192 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 23109 20791 23167 20797
rect 23109 20788 23121 20791
rect 22888 20760 23121 20788
rect 22888 20748 22894 20760
rect 23109 20757 23121 20760
rect 23155 20757 23167 20791
rect 23216 20788 23244 20896
rect 23293 20893 23305 20927
rect 23339 20924 23351 20927
rect 23474 20924 23480 20936
rect 23339 20896 23480 20924
rect 23339 20893 23351 20896
rect 23293 20887 23351 20893
rect 23474 20884 23480 20896
rect 23532 20884 23538 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 25314 20924 25320 20936
rect 23615 20896 25320 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20924 25467 20927
rect 26786 20924 26792 20936
rect 25455 20896 26792 20924
rect 25455 20893 25467 20896
rect 25409 20887 25467 20893
rect 26786 20884 26792 20896
rect 26844 20924 26850 20936
rect 27430 20924 27436 20936
rect 26844 20896 27436 20924
rect 26844 20884 26850 20896
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27522 20884 27528 20936
rect 27580 20924 27586 20936
rect 28843 20933 28871 20964
rect 29086 20952 29092 21004
rect 29144 20992 29150 21004
rect 30760 21001 30788 21032
rect 31021 21029 31033 21063
rect 31067 21060 31079 21063
rect 32677 21063 32735 21069
rect 31067 21032 32444 21060
rect 31067 21029 31079 21032
rect 31021 21023 31079 21029
rect 29825 20995 29883 21001
rect 29825 20992 29837 20995
rect 29144 20964 29837 20992
rect 29144 20952 29150 20964
rect 29825 20961 29837 20964
rect 29871 20961 29883 20995
rect 29825 20955 29883 20961
rect 30745 20995 30803 21001
rect 30745 20961 30757 20995
rect 30791 20961 30803 20995
rect 30745 20955 30803 20961
rect 28537 20927 28595 20933
rect 27580 20896 27625 20924
rect 27580 20884 27586 20896
rect 28537 20893 28549 20927
rect 28583 20893 28595 20927
rect 28631 20927 28689 20933
rect 28631 20914 28643 20927
rect 28677 20914 28689 20927
rect 28843 20927 28917 20933
rect 28537 20887 28595 20893
rect 24210 20816 24216 20868
rect 24268 20856 24274 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 24268 20828 24593 20856
rect 24268 20816 24274 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24581 20819 24639 20825
rect 24797 20859 24855 20865
rect 24797 20825 24809 20859
rect 24843 20856 24855 20859
rect 25498 20856 25504 20868
rect 24843 20828 25504 20856
rect 24843 20825 24855 20828
rect 24797 20819 24855 20825
rect 25498 20816 25504 20828
rect 25556 20816 25562 20868
rect 25676 20859 25734 20865
rect 25676 20825 25688 20859
rect 25722 20856 25734 20859
rect 26234 20856 26240 20868
rect 25722 20828 26240 20856
rect 25722 20825 25734 20828
rect 25676 20819 25734 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 27801 20859 27859 20865
rect 27801 20825 27813 20859
rect 27847 20825 27859 20859
rect 27801 20819 27859 20825
rect 23566 20788 23572 20800
rect 23216 20760 23572 20788
rect 23109 20751 23167 20757
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 26418 20788 26424 20800
rect 24995 20760 26424 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 27816 20788 27844 20819
rect 28442 20816 28448 20868
rect 28500 20856 28506 20868
rect 28552 20856 28580 20887
rect 28626 20862 28632 20914
rect 28684 20862 28690 20914
rect 28843 20896 28871 20927
rect 28859 20893 28871 20896
rect 28905 20893 28917 20927
rect 28994 20924 29000 20936
rect 28955 20896 29000 20924
rect 28859 20887 28917 20893
rect 28994 20884 29000 20896
rect 29052 20924 29058 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29052 20896 29745 20924
rect 29052 20884 29058 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 30193 20927 30251 20933
rect 30193 20893 30205 20927
rect 30239 20893 30251 20927
rect 30193 20887 30251 20893
rect 28500 20828 28580 20856
rect 28500 20816 28506 20828
rect 28718 20816 28724 20868
rect 28776 20856 28782 20868
rect 29086 20856 29092 20868
rect 28776 20828 29092 20856
rect 28776 20816 28782 20828
rect 29086 20816 29092 20828
rect 29144 20816 29150 20868
rect 29178 20816 29184 20868
rect 29236 20856 29242 20868
rect 30208 20856 30236 20887
rect 30558 20884 30564 20936
rect 30616 20924 30622 20936
rect 31588 20933 31616 21032
rect 32416 21004 32444 21032
rect 32677 21029 32689 21063
rect 32723 21060 32735 21063
rect 32766 21060 32772 21072
rect 32723 21032 32772 21060
rect 32723 21029 32735 21032
rect 32677 21023 32735 21029
rect 32766 21020 32772 21032
rect 32824 21020 32830 21072
rect 32858 21020 32864 21072
rect 32916 21060 32922 21072
rect 32916 21032 34008 21060
rect 32916 21020 32922 21032
rect 31849 20995 31907 21001
rect 31849 20961 31861 20995
rect 31895 20992 31907 20995
rect 31895 20964 32352 20992
rect 31895 20961 31907 20964
rect 31849 20955 31907 20961
rect 32324 20936 32352 20964
rect 32398 20952 32404 21004
rect 32456 20992 32462 21004
rect 32456 20964 33272 20992
rect 32456 20952 32462 20964
rect 30653 20927 30711 20933
rect 30653 20924 30665 20927
rect 30616 20896 30665 20924
rect 30616 20884 30622 20896
rect 30653 20893 30665 20896
rect 30699 20893 30711 20927
rect 30653 20887 30711 20893
rect 31573 20927 31631 20933
rect 31573 20893 31585 20927
rect 31619 20893 31631 20927
rect 32306 20924 32312 20936
rect 32267 20896 32312 20924
rect 31573 20887 31631 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 33137 20927 33195 20933
rect 33137 20893 33149 20927
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 29236 20828 30236 20856
rect 31849 20859 31907 20865
rect 29236 20816 29242 20828
rect 31849 20825 31861 20859
rect 31895 20856 31907 20859
rect 33152 20856 33180 20887
rect 31895 20828 33180 20856
rect 33244 20856 33272 20964
rect 33318 20952 33324 21004
rect 33376 20992 33382 21004
rect 33376 20964 33421 20992
rect 33376 20952 33382 20964
rect 33505 20927 33563 20933
rect 33505 20893 33517 20927
rect 33551 20918 33563 20927
rect 33870 20924 33876 20936
rect 33612 20918 33876 20924
rect 33551 20896 33876 20918
rect 33551 20893 33640 20896
rect 33505 20890 33640 20893
rect 33505 20887 33563 20890
rect 33870 20884 33876 20896
rect 33928 20884 33934 20936
rect 33980 20933 34008 21032
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20893 34207 20927
rect 34149 20887 34207 20893
rect 34164 20856 34192 20887
rect 33244 20828 34192 20856
rect 31895 20825 31907 20828
rect 31849 20819 31907 20825
rect 29546 20788 29552 20800
rect 27816 20760 29552 20788
rect 29546 20748 29552 20760
rect 29604 20748 29610 20800
rect 29822 20748 29828 20800
rect 29880 20788 29886 20800
rect 29917 20791 29975 20797
rect 29917 20788 29929 20791
rect 29880 20760 29929 20788
rect 29880 20748 29886 20760
rect 29917 20757 29929 20760
rect 29963 20757 29975 20791
rect 29917 20751 29975 20757
rect 30101 20791 30159 20797
rect 30101 20757 30113 20791
rect 30147 20788 30159 20791
rect 30834 20788 30840 20800
rect 30147 20760 30840 20788
rect 30147 20757 30159 20760
rect 30101 20751 30159 20757
rect 30834 20748 30840 20760
rect 30892 20748 30898 20800
rect 32766 20748 32772 20800
rect 32824 20788 32830 20800
rect 33229 20791 33287 20797
rect 33229 20788 33241 20791
rect 32824 20760 33241 20788
rect 32824 20748 32830 20760
rect 33229 20757 33241 20760
rect 33275 20757 33287 20791
rect 33410 20788 33416 20800
rect 33371 20760 33416 20788
rect 33229 20751 33287 20757
rect 33410 20748 33416 20760
rect 33468 20748 33474 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12860 20556 12909 20584
rect 12860 20544 12866 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 15013 20587 15071 20593
rect 15013 20553 15025 20587
rect 15059 20584 15071 20587
rect 15102 20584 15108 20596
rect 15059 20556 15108 20584
rect 15059 20553 15071 20556
rect 15013 20547 15071 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 19981 20587 20039 20593
rect 19981 20584 19993 20587
rect 18564 20556 19993 20584
rect 18564 20544 18570 20556
rect 19981 20553 19993 20556
rect 20027 20553 20039 20587
rect 19981 20547 20039 20553
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 21692 20556 22048 20584
rect 21692 20544 21698 20556
rect 13446 20476 13452 20528
rect 13504 20516 13510 20528
rect 15933 20519 15991 20525
rect 15933 20516 15945 20519
rect 13504 20488 15945 20516
rect 13504 20476 13510 20488
rect 15933 20485 15945 20488
rect 15979 20485 15991 20519
rect 15933 20479 15991 20485
rect 18046 20476 18052 20528
rect 18104 20516 18110 20528
rect 18202 20519 18260 20525
rect 18202 20516 18214 20519
rect 18104 20488 18214 20516
rect 18104 20476 18110 20488
rect 18202 20485 18214 20488
rect 18248 20485 18260 20519
rect 18202 20479 18260 20485
rect 20901 20519 20959 20525
rect 20901 20485 20913 20519
rect 20947 20516 20959 20519
rect 20990 20516 20996 20528
rect 20947 20488 20996 20516
rect 20947 20485 20959 20488
rect 20901 20479 20959 20485
rect 20990 20476 20996 20488
rect 21048 20476 21054 20528
rect 22020 20525 22048 20556
rect 22646 20544 22652 20596
rect 22704 20584 22710 20596
rect 23198 20584 23204 20596
rect 22704 20556 23204 20584
rect 22704 20544 22710 20556
rect 23198 20544 23204 20556
rect 23256 20544 23262 20596
rect 26234 20584 26240 20596
rect 26195 20556 26240 20584
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 26418 20544 26424 20596
rect 26476 20544 26482 20596
rect 28445 20587 28503 20593
rect 28445 20553 28457 20587
rect 28491 20584 28503 20587
rect 28534 20584 28540 20596
rect 28491 20556 28540 20584
rect 28491 20553 28503 20556
rect 28445 20547 28503 20553
rect 28534 20544 28540 20556
rect 28592 20544 28598 20596
rect 28626 20544 28632 20596
rect 28684 20584 28690 20596
rect 28902 20584 28908 20596
rect 28684 20556 28908 20584
rect 28684 20544 28690 20556
rect 28902 20544 28908 20556
rect 28960 20584 28966 20596
rect 29822 20584 29828 20596
rect 28960 20556 29828 20584
rect 28960 20544 28966 20556
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 32309 20587 32367 20593
rect 32309 20553 32321 20587
rect 32355 20584 32367 20587
rect 32582 20584 32588 20596
rect 32355 20556 32588 20584
rect 32355 20553 32367 20556
rect 32309 20547 32367 20553
rect 32582 20544 32588 20556
rect 32640 20544 32646 20596
rect 32677 20587 32735 20593
rect 32677 20553 32689 20587
rect 32723 20584 32735 20587
rect 32766 20584 32772 20596
rect 32723 20556 32772 20584
rect 32723 20553 32735 20556
rect 32677 20547 32735 20553
rect 32766 20544 32772 20556
rect 32824 20584 32830 20596
rect 32950 20584 32956 20596
rect 32824 20556 32956 20584
rect 32824 20544 32830 20556
rect 32950 20544 32956 20556
rect 33008 20544 33014 20596
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 34885 20587 34943 20593
rect 34885 20584 34897 20587
rect 34848 20556 34897 20584
rect 34848 20544 34854 20556
rect 34885 20553 34897 20556
rect 34931 20553 34943 20587
rect 34885 20547 34943 20553
rect 22005 20519 22063 20525
rect 22005 20485 22017 20519
rect 22051 20485 22063 20519
rect 22005 20479 22063 20485
rect 12618 20408 12624 20460
rect 12676 20448 12682 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12676 20420 12817 20448
rect 12676 20408 12682 20420
rect 12805 20417 12817 20420
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20448 13691 20451
rect 13722 20448 13728 20460
rect 13679 20420 13728 20448
rect 13679 20417 13691 20420
rect 13633 20411 13691 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 13906 20457 13912 20460
rect 13900 20411 13912 20457
rect 13964 20448 13970 20460
rect 13964 20420 14000 20448
rect 13906 20408 13912 20411
rect 13964 20408 13970 20420
rect 16390 20408 16396 20460
rect 16448 20448 16454 20460
rect 17957 20451 18015 20457
rect 17957 20448 17969 20451
rect 16448 20420 17969 20448
rect 16448 20408 16454 20420
rect 17957 20417 17969 20420
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 19242 20408 19248 20460
rect 19300 20448 19306 20460
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 19300 20420 19901 20448
rect 19300 20408 19306 20420
rect 19889 20417 19901 20420
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 21082 20408 21088 20460
rect 21140 20448 21146 20460
rect 21634 20448 21640 20460
rect 21140 20420 21640 20448
rect 21140 20408 21146 20420
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 21726 20408 21732 20460
rect 21784 20448 21790 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21784 20420 21833 20448
rect 21784 20408 21790 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 23106 20448 23112 20460
rect 23067 20420 23112 20448
rect 21821 20411 21879 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23382 20457 23388 20460
rect 23376 20411 23388 20457
rect 23440 20448 23446 20460
rect 23440 20420 23476 20448
rect 23382 20408 23388 20411
rect 23440 20408 23446 20420
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 26436 20457 26464 20544
rect 27246 20476 27252 20528
rect 27304 20516 27310 20528
rect 27304 20488 27476 20516
rect 27304 20476 27310 20488
rect 27448 20457 27476 20488
rect 33410 20476 33416 20528
rect 33468 20516 33474 20528
rect 33750 20519 33808 20525
rect 33750 20516 33762 20519
rect 33468 20488 33762 20516
rect 33468 20476 33474 20488
rect 33750 20485 33762 20488
rect 33796 20485 33808 20519
rect 33750 20479 33808 20485
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24912 20420 24961 20448
rect 24912 20408 24918 20420
rect 24949 20417 24961 20420
rect 24995 20417 25007 20451
rect 24949 20411 25007 20417
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20417 26479 20451
rect 26421 20411 26479 20417
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 15470 20340 15476 20392
rect 15528 20380 15534 20392
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 15528 20352 16681 20380
rect 15528 20340 15534 20352
rect 16669 20349 16681 20352
rect 16715 20349 16727 20383
rect 16942 20380 16948 20392
rect 16903 20352 16948 20380
rect 16669 20343 16727 20349
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 20438 20340 20444 20392
rect 20496 20380 20502 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20496 20352 21005 20380
rect 20496 20340 20502 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 21174 20380 21180 20392
rect 21135 20352 21180 20380
rect 20993 20343 21051 20349
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 24670 20340 24676 20392
rect 24728 20380 24734 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 24728 20352 25237 20380
rect 24728 20340 24734 20352
rect 25225 20349 25237 20352
rect 25271 20349 25283 20383
rect 25225 20343 25283 20349
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 25556 20352 26985 20380
rect 25556 20340 25562 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 27157 20383 27215 20389
rect 27157 20349 27169 20383
rect 27203 20349 27215 20383
rect 27157 20343 27215 20349
rect 27249 20383 27307 20389
rect 27249 20349 27261 20383
rect 27295 20349 27307 20383
rect 27356 20380 27384 20411
rect 27798 20408 27804 20460
rect 27856 20448 27862 20460
rect 28629 20451 28687 20457
rect 28629 20448 28641 20451
rect 27856 20420 28641 20448
rect 27856 20408 27862 20420
rect 28629 20417 28641 20420
rect 28675 20417 28687 20451
rect 28629 20411 28687 20417
rect 28997 20451 29055 20457
rect 28997 20417 29009 20451
rect 29043 20448 29055 20451
rect 29730 20448 29736 20460
rect 29043 20420 29736 20448
rect 29043 20417 29055 20420
rect 28997 20411 29055 20417
rect 29730 20408 29736 20420
rect 29788 20408 29794 20460
rect 30282 20448 30288 20460
rect 30243 20420 30288 20448
rect 30282 20408 30288 20420
rect 30340 20408 30346 20460
rect 31386 20448 31392 20460
rect 31347 20420 31392 20448
rect 31386 20408 31392 20420
rect 31444 20408 31450 20460
rect 32769 20451 32827 20457
rect 32769 20417 32781 20451
rect 32815 20448 32827 20451
rect 33318 20448 33324 20460
rect 32815 20420 33324 20448
rect 32815 20417 32827 20420
rect 32769 20411 32827 20417
rect 33318 20408 33324 20420
rect 33376 20408 33382 20460
rect 33502 20448 33508 20460
rect 33463 20420 33508 20448
rect 33502 20408 33508 20420
rect 33560 20408 33566 20460
rect 27356 20352 27476 20380
rect 27249 20343 27307 20349
rect 19058 20272 19064 20324
rect 19116 20312 19122 20324
rect 19337 20315 19395 20321
rect 19337 20312 19349 20315
rect 19116 20284 19349 20312
rect 19116 20272 19122 20284
rect 19337 20281 19349 20284
rect 19383 20312 19395 20315
rect 20456 20312 20484 20340
rect 19383 20284 20484 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 25590 20272 25596 20324
rect 25648 20312 25654 20324
rect 27172 20312 27200 20343
rect 25648 20284 27200 20312
rect 27264 20312 27292 20343
rect 27338 20312 27344 20324
rect 27264 20284 27344 20312
rect 25648 20272 25654 20284
rect 27338 20272 27344 20284
rect 27396 20272 27402 20324
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15620 20216 16037 20244
rect 15620 20204 15626 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 20533 20247 20591 20253
rect 20533 20213 20545 20247
rect 20579 20244 20591 20247
rect 21174 20244 21180 20256
rect 20579 20216 21180 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 22189 20247 22247 20253
rect 22189 20213 22201 20247
rect 22235 20244 22247 20247
rect 23106 20244 23112 20256
rect 22235 20216 23112 20244
rect 22235 20213 22247 20216
rect 22189 20207 22247 20213
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24489 20247 24547 20253
rect 24489 20244 24501 20247
rect 24360 20216 24501 20244
rect 24360 20204 24366 20216
rect 24489 20213 24501 20216
rect 24535 20244 24547 20247
rect 27448 20244 27476 20352
rect 28534 20340 28540 20392
rect 28592 20380 28598 20392
rect 28718 20380 28724 20392
rect 28592 20352 28724 20380
rect 28592 20340 28598 20352
rect 28718 20340 28724 20352
rect 28776 20340 28782 20392
rect 29089 20383 29147 20389
rect 29089 20349 29101 20383
rect 29135 20349 29147 20383
rect 30377 20383 30435 20389
rect 30377 20380 30389 20383
rect 29089 20343 29147 20349
rect 30300 20352 30389 20380
rect 28074 20272 28080 20324
rect 28132 20312 28138 20324
rect 29104 20312 29132 20343
rect 30300 20324 30328 20352
rect 30377 20349 30389 20352
rect 30423 20349 30435 20383
rect 30377 20343 30435 20349
rect 30466 20340 30472 20392
rect 30524 20380 30530 20392
rect 32861 20383 32919 20389
rect 32861 20380 32873 20383
rect 30524 20352 30569 20380
rect 31726 20352 32873 20380
rect 30524 20340 30530 20352
rect 29914 20312 29920 20324
rect 28132 20284 29132 20312
rect 29875 20284 29920 20312
rect 28132 20272 28138 20284
rect 24535 20216 27476 20244
rect 24535 20213 24547 20216
rect 24489 20207 24547 20213
rect 28166 20204 28172 20256
rect 28224 20244 28230 20256
rect 28718 20244 28724 20256
rect 28224 20216 28724 20244
rect 28224 20204 28230 20216
rect 28718 20204 28724 20216
rect 28776 20204 28782 20256
rect 29104 20244 29132 20284
rect 29914 20272 29920 20284
rect 29972 20272 29978 20324
rect 30282 20272 30288 20324
rect 30340 20272 30346 20324
rect 31481 20247 31539 20253
rect 31481 20244 31493 20247
rect 29104 20216 31493 20244
rect 31481 20213 31493 20216
rect 31527 20244 31539 20247
rect 31726 20244 31754 20352
rect 32861 20349 32873 20352
rect 32907 20349 32919 20383
rect 32861 20343 32919 20349
rect 31527 20216 31754 20244
rect 31527 20213 31539 20216
rect 31481 20207 31539 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13906 20040 13912 20052
rect 13403 20012 13912 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 19797 20043 19855 20049
rect 19797 20009 19809 20043
rect 19843 20040 19855 20043
rect 20530 20040 20536 20052
rect 19843 20012 20536 20040
rect 19843 20009 19855 20012
rect 19797 20003 19855 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 20916 20012 21404 20040
rect 17310 19932 17316 19984
rect 17368 19972 17374 19984
rect 17368 19944 18092 19972
rect 17368 19932 17374 19944
rect 15378 19904 15384 19916
rect 14292 19876 15384 19904
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 13541 19799 13599 19805
rect 13556 19768 13584 19799
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14292 19845 14320 19876
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 17034 19864 17040 19916
rect 17092 19904 17098 19916
rect 17862 19904 17868 19916
rect 17092 19876 17868 19904
rect 17092 19864 17098 19876
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 15013 19839 15071 19845
rect 15013 19805 15025 19839
rect 15059 19836 15071 19839
rect 15562 19836 15568 19848
rect 15059 19808 15568 19836
rect 15059 19805 15071 19808
rect 15013 19799 15071 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 16206 19836 16212 19848
rect 15703 19808 16212 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 14461 19771 14519 19777
rect 14461 19768 14473 19771
rect 13556 19740 14473 19768
rect 14461 19737 14473 19740
rect 14507 19737 14519 19771
rect 14461 19731 14519 19737
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15672 19768 15700 19799
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17497 19839 17555 19845
rect 17497 19836 17509 19839
rect 17000 19808 17509 19836
rect 17000 19796 17006 19808
rect 17497 19805 17509 19808
rect 17543 19805 17555 19839
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17497 19799 17555 19805
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 18064 19845 18092 19944
rect 20714 19932 20720 19984
rect 20772 19972 20778 19984
rect 20809 19975 20867 19981
rect 20809 19972 20821 19975
rect 20772 19944 20821 19972
rect 20772 19932 20778 19944
rect 20809 19941 20821 19944
rect 20855 19941 20867 19975
rect 20809 19935 20867 19941
rect 20165 19907 20223 19913
rect 20165 19873 20177 19907
rect 20211 19904 20223 19907
rect 20916 19904 20944 20012
rect 20211 19876 20944 19904
rect 21376 19904 21404 20012
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 21913 20043 21971 20049
rect 21913 20040 21925 20043
rect 21508 20012 21925 20040
rect 21508 20000 21514 20012
rect 21913 20009 21925 20012
rect 21959 20009 21971 20043
rect 23382 20040 23388 20052
rect 23343 20012 23388 20040
rect 21913 20003 21971 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 24578 20040 24584 20052
rect 24412 20012 24584 20040
rect 22094 19932 22100 19984
rect 22152 19932 22158 19984
rect 22186 19932 22192 19984
rect 22244 19972 22250 19984
rect 23753 19975 23811 19981
rect 23753 19972 23765 19975
rect 22244 19944 23765 19972
rect 22244 19932 22250 19944
rect 23753 19941 23765 19944
rect 23799 19941 23811 19975
rect 23753 19935 23811 19941
rect 22112 19904 22140 19932
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 21376 19876 22293 19904
rect 20211 19873 20223 19876
rect 20165 19867 20223 19873
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 24412 19904 24440 20012
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 26329 20043 26387 20049
rect 26329 20009 26341 20043
rect 26375 20040 26387 20043
rect 27522 20040 27528 20052
rect 26375 20012 27528 20040
rect 26375 20009 26387 20012
rect 26329 20003 26387 20009
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 27709 20043 27767 20049
rect 27709 20009 27721 20043
rect 27755 20040 27767 20043
rect 30558 20040 30564 20052
rect 27755 20012 29776 20040
rect 30519 20012 30564 20040
rect 27755 20009 27767 20012
rect 27709 20003 27767 20009
rect 24486 19932 24492 19984
rect 24544 19972 24550 19984
rect 24857 19975 24915 19981
rect 24544 19944 24808 19972
rect 24544 19932 24550 19944
rect 24780 19904 24808 19944
rect 24857 19941 24869 19975
rect 24903 19972 24915 19975
rect 25130 19972 25136 19984
rect 24903 19944 25136 19972
rect 24903 19941 24915 19944
rect 24857 19935 24915 19941
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 27617 19975 27675 19981
rect 27617 19941 27629 19975
rect 27663 19972 27675 19975
rect 28074 19972 28080 19984
rect 27663 19944 28080 19972
rect 27663 19941 27675 19944
rect 27617 19935 27675 19941
rect 28074 19932 28080 19944
rect 28132 19932 28138 19984
rect 29748 19972 29776 20012
rect 30558 20000 30564 20012
rect 30616 20000 30622 20052
rect 32401 20043 32459 20049
rect 32401 20009 32413 20043
rect 32447 20040 32459 20043
rect 32858 20040 32864 20052
rect 32447 20012 32864 20040
rect 32447 20009 32459 20012
rect 32401 20003 32459 20009
rect 32858 20000 32864 20012
rect 32916 20000 32922 20052
rect 35342 19972 35348 19984
rect 29748 19944 35204 19972
rect 35303 19944 35348 19972
rect 28445 19907 28503 19913
rect 28445 19904 28457 19907
rect 24412 19876 24716 19904
rect 24780 19876 28457 19904
rect 22281 19867 22339 19873
rect 18049 19839 18107 19845
rect 17828 19808 17873 19836
rect 17828 19796 17834 19808
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 19978 19836 19984 19848
rect 19939 19808 19984 19836
rect 18049 19799 18107 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19805 20131 19839
rect 20254 19836 20260 19848
rect 20215 19808 20260 19836
rect 20073 19799 20131 19805
rect 15243 19740 15700 19768
rect 15924 19771 15982 19777
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15924 19737 15936 19771
rect 15970 19768 15982 19771
rect 16390 19768 16396 19780
rect 15970 19740 16396 19768
rect 15970 19737 15982 19740
rect 15924 19731 15982 19737
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 18782 19768 18788 19780
rect 17052 19740 18788 19768
rect 16942 19660 16948 19712
rect 17000 19700 17006 19712
rect 17052 19709 17080 19740
rect 18782 19728 18788 19740
rect 18840 19728 18846 19780
rect 20088 19768 20116 19799
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 20622 19796 20628 19848
rect 20680 19836 20686 19848
rect 21085 19839 21143 19845
rect 21290 19839 21348 19845
rect 21085 19838 21097 19839
rect 21080 19836 21097 19838
rect 20680 19808 21097 19836
rect 20680 19796 20686 19808
rect 21054 19805 21097 19808
rect 21131 19805 21143 19839
rect 21054 19802 21143 19805
rect 21085 19799 21143 19802
rect 21190 19833 21248 19839
rect 21190 19799 21202 19833
rect 21236 19799 21248 19833
rect 21290 19805 21302 19839
rect 21336 19836 21348 19839
rect 21336 19808 21404 19836
rect 21336 19805 21348 19808
rect 21290 19799 21348 19805
rect 21190 19793 21248 19799
rect 20714 19768 20720 19780
rect 20088 19740 20720 19768
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 21192 19712 21220 19793
rect 17037 19703 17095 19709
rect 17037 19700 17049 19703
rect 17000 19672 17049 19700
rect 17000 19660 17006 19672
rect 17037 19669 17049 19672
rect 17083 19669 17095 19703
rect 17037 19663 17095 19669
rect 18233 19703 18291 19709
rect 18233 19669 18245 19703
rect 18279 19700 18291 19703
rect 18322 19700 18328 19712
rect 18279 19672 18328 19700
rect 18279 19669 18291 19672
rect 18233 19663 18291 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 21174 19660 21180 19712
rect 21232 19660 21238 19712
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21376 19700 21404 19808
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 22094 19836 22100 19848
rect 21508 19808 21553 19836
rect 22055 19808 22100 19836
rect 21508 19796 21514 19808
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22244 19808 22289 19836
rect 22244 19796 22250 19808
rect 22370 19796 22376 19848
rect 22428 19836 22434 19848
rect 22428 19808 22473 19836
rect 22428 19796 22434 19808
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23532 19808 23581 19836
rect 23532 19796 23538 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19836 23903 19839
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23891 19808 24593 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24688 19836 24716 19876
rect 28445 19873 28457 19876
rect 28491 19873 28503 19907
rect 31113 19907 31171 19913
rect 31113 19904 31125 19907
rect 28445 19867 28503 19873
rect 30576 19876 31125 19904
rect 24765 19839 24823 19845
rect 24765 19836 24777 19839
rect 24688 19808 24777 19836
rect 24581 19799 24639 19805
rect 24765 19805 24777 19808
rect 24811 19805 24823 19839
rect 24765 19799 24823 19805
rect 23584 19768 23612 19799
rect 24854 19796 24860 19848
rect 24912 19836 24918 19848
rect 24949 19839 25007 19845
rect 24949 19836 24961 19839
rect 24912 19808 24961 19836
rect 24912 19796 24918 19808
rect 24949 19805 24961 19808
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 24670 19768 24676 19780
rect 23584 19740 24676 19768
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 25056 19768 25084 19799
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25961 19839 26019 19845
rect 25961 19836 25973 19839
rect 25832 19808 25973 19836
rect 25832 19796 25838 19808
rect 25961 19805 25973 19808
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19836 26387 19839
rect 26510 19836 26516 19848
rect 26375 19808 26516 19836
rect 26375 19805 26387 19808
rect 26329 19799 26387 19805
rect 26510 19796 26516 19808
rect 26568 19796 26574 19848
rect 29546 19796 29552 19848
rect 29604 19836 29610 19848
rect 29917 19839 29975 19845
rect 29917 19836 29929 19839
rect 29604 19808 29929 19836
rect 29604 19796 29610 19808
rect 29917 19805 29929 19808
rect 29963 19836 29975 19839
rect 30466 19836 30472 19848
rect 29963 19808 30472 19836
rect 29963 19805 29975 19808
rect 29917 19799 29975 19805
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 27246 19768 27252 19780
rect 24964 19740 25084 19768
rect 27207 19740 27252 19768
rect 21324 19672 21404 19700
rect 21324 19660 21330 19672
rect 21450 19660 21456 19712
rect 21508 19700 21514 19712
rect 21818 19700 21824 19712
rect 21508 19672 21824 19700
rect 21508 19660 21514 19672
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 24302 19700 24308 19712
rect 23532 19672 24308 19700
rect 23532 19660 23538 19672
rect 24302 19660 24308 19672
rect 24360 19700 24366 19712
rect 24964 19700 24992 19740
rect 27246 19728 27252 19740
rect 27304 19728 27310 19780
rect 28258 19768 28264 19780
rect 28219 19740 28264 19768
rect 28258 19728 28264 19740
rect 28316 19768 28322 19780
rect 28810 19768 28816 19780
rect 28316 19740 28816 19768
rect 28316 19728 28322 19740
rect 28810 19728 28816 19740
rect 28868 19728 28874 19780
rect 30576 19768 30604 19876
rect 31113 19873 31125 19876
rect 31159 19904 31171 19907
rect 31386 19904 31392 19916
rect 31159 19876 31392 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 31386 19864 31392 19876
rect 31444 19904 31450 19916
rect 32953 19907 33011 19913
rect 32953 19904 32965 19907
rect 31444 19876 32965 19904
rect 31444 19864 31450 19876
rect 32953 19873 32965 19876
rect 32999 19904 33011 19907
rect 33134 19904 33140 19916
rect 32999 19876 33140 19904
rect 32999 19873 33011 19876
rect 32953 19867 33011 19873
rect 33134 19864 33140 19876
rect 33192 19864 33198 19916
rect 30650 19796 30656 19848
rect 30708 19836 30714 19848
rect 30926 19836 30932 19848
rect 30708 19808 30932 19836
rect 30708 19796 30714 19808
rect 30926 19796 30932 19808
rect 30984 19796 30990 19848
rect 31018 19796 31024 19848
rect 31076 19836 31082 19848
rect 31757 19839 31815 19845
rect 31757 19836 31769 19839
rect 31076 19808 31769 19836
rect 31076 19796 31082 19808
rect 31757 19805 31769 19808
rect 31803 19805 31815 19839
rect 31757 19799 31815 19805
rect 32582 19796 32588 19848
rect 32640 19836 32646 19848
rect 32769 19839 32827 19845
rect 32769 19836 32781 19839
rect 32640 19808 32781 19836
rect 32640 19796 32646 19808
rect 32769 19805 32781 19808
rect 32815 19836 32827 19839
rect 33042 19836 33048 19848
rect 32815 19808 33048 19836
rect 32815 19805 32827 19808
rect 32769 19799 32827 19805
rect 33042 19796 33048 19808
rect 33100 19796 33106 19848
rect 33410 19796 33416 19848
rect 33468 19836 33474 19848
rect 35176 19845 35204 19944
rect 35342 19932 35348 19944
rect 35400 19932 35406 19984
rect 33597 19839 33655 19845
rect 33597 19836 33609 19839
rect 33468 19808 33609 19836
rect 33468 19796 33474 19808
rect 33597 19805 33609 19808
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 35161 19839 35219 19845
rect 35161 19805 35173 19839
rect 35207 19805 35219 19839
rect 35161 19799 35219 19805
rect 30024 19740 30604 19768
rect 32861 19771 32919 19777
rect 24360 19672 24992 19700
rect 24360 19660 24366 19672
rect 25314 19660 25320 19712
rect 25372 19700 25378 19712
rect 26513 19703 26571 19709
rect 26513 19700 26525 19703
rect 25372 19672 26525 19700
rect 25372 19660 25378 19672
rect 26513 19669 26525 19672
rect 26559 19669 26571 19703
rect 26513 19663 26571 19669
rect 28442 19660 28448 19712
rect 28500 19700 28506 19712
rect 30024 19709 30052 19740
rect 32861 19737 32873 19771
rect 32907 19768 32919 19771
rect 33778 19768 33784 19780
rect 32907 19740 33784 19768
rect 32907 19737 32919 19740
rect 32861 19731 32919 19737
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 30009 19703 30067 19709
rect 30009 19700 30021 19703
rect 28500 19672 30021 19700
rect 28500 19660 28506 19672
rect 30009 19669 30021 19672
rect 30055 19669 30067 19703
rect 30009 19663 30067 19669
rect 31021 19703 31079 19709
rect 31021 19669 31033 19703
rect 31067 19700 31079 19703
rect 31849 19703 31907 19709
rect 31849 19700 31861 19703
rect 31067 19672 31861 19700
rect 31067 19669 31079 19672
rect 31021 19663 31079 19669
rect 31849 19669 31861 19672
rect 31895 19669 31907 19703
rect 31849 19663 31907 19669
rect 32950 19660 32956 19712
rect 33008 19700 33014 19712
rect 33689 19703 33747 19709
rect 33689 19700 33701 19703
rect 33008 19672 33701 19700
rect 33008 19660 33014 19672
rect 33689 19669 33701 19672
rect 33735 19669 33747 19703
rect 33689 19663 33747 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 19429 19499 19487 19505
rect 19429 19465 19441 19499
rect 19475 19496 19487 19499
rect 20254 19496 20260 19508
rect 19475 19468 20260 19496
rect 19475 19465 19487 19468
rect 19429 19459 19487 19465
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20364 19468 20944 19496
rect 13446 19428 13452 19440
rect 13407 19400 13452 19428
rect 13446 19388 13452 19400
rect 13504 19388 13510 19440
rect 14737 19431 14795 19437
rect 14737 19397 14749 19431
rect 14783 19428 14795 19431
rect 17126 19428 17132 19440
rect 14783 19400 17132 19428
rect 14783 19397 14795 19400
rect 14737 19391 14795 19397
rect 17126 19388 17132 19400
rect 17184 19428 17190 19440
rect 19242 19428 19248 19440
rect 17184 19400 19248 19428
rect 17184 19388 17190 19400
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 20364 19428 20392 19468
rect 20916 19437 20944 19468
rect 20990 19456 20996 19508
rect 21048 19456 21054 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 22186 19496 22192 19508
rect 21223 19468 22192 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 24765 19499 24823 19505
rect 24765 19465 24777 19499
rect 24811 19496 24823 19499
rect 25038 19496 25044 19508
rect 24811 19468 25044 19496
rect 24811 19465 24823 19468
rect 24765 19459 24823 19465
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 26973 19499 27031 19505
rect 26973 19465 26985 19499
rect 27019 19496 27031 19499
rect 27246 19496 27252 19508
rect 27019 19468 27252 19496
rect 27019 19465 27031 19468
rect 26973 19459 27031 19465
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 27430 19496 27436 19508
rect 27391 19468 27436 19496
rect 27430 19456 27436 19468
rect 27488 19456 27494 19508
rect 28074 19496 28080 19508
rect 28035 19468 28080 19496
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 32306 19456 32312 19508
rect 32364 19496 32370 19508
rect 32493 19499 32551 19505
rect 32493 19496 32505 19499
rect 32364 19468 32505 19496
rect 32364 19456 32370 19468
rect 32493 19465 32505 19468
rect 32539 19465 32551 19499
rect 32950 19496 32956 19508
rect 32911 19468 32956 19496
rect 32493 19459 32551 19465
rect 32950 19456 32956 19468
rect 33008 19456 33014 19508
rect 33778 19496 33784 19508
rect 33739 19468 33784 19496
rect 33778 19456 33784 19468
rect 33836 19456 33842 19508
rect 19352 19400 20392 19428
rect 20901 19431 20959 19437
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12253 19363 12311 19369
rect 12253 19360 12265 19363
rect 11940 19332 12265 19360
rect 11940 19320 11946 19332
rect 12253 19329 12265 19332
rect 12299 19329 12311 19363
rect 12253 19323 12311 19329
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 15436 19332 15485 19360
rect 15436 19320 15442 19332
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16850 19360 16856 19372
rect 16811 19332 16856 19360
rect 16669 19323 16727 19329
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15102 19224 15108 19236
rect 14967 19196 15108 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15102 19184 15108 19196
rect 15160 19184 15166 19236
rect 16684 19224 16712 19323
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 17034 19360 17040 19372
rect 16995 19332 17040 19360
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17218 19360 17224 19372
rect 17179 19332 17224 19360
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 18322 19360 18328 19372
rect 18283 19332 18328 19360
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18506 19360 18512 19372
rect 18467 19332 18512 19360
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 19352 19360 19380 19400
rect 20901 19397 20913 19431
rect 20947 19397 20959 19431
rect 21008 19428 21036 19456
rect 21818 19428 21824 19440
rect 21008 19400 21824 19428
rect 20901 19391 20959 19397
rect 21818 19388 21824 19400
rect 21876 19388 21882 19440
rect 21913 19431 21971 19437
rect 21913 19397 21925 19431
rect 21959 19428 21971 19431
rect 24486 19428 24492 19440
rect 21959 19400 24492 19428
rect 21959 19397 21971 19400
rect 21913 19391 21971 19397
rect 24486 19388 24492 19400
rect 24544 19388 24550 19440
rect 27448 19428 27476 19456
rect 24780 19400 26234 19428
rect 27448 19400 28580 19428
rect 24780 19372 24808 19400
rect 18840 19332 19380 19360
rect 19705 19363 19763 19369
rect 18840 19320 18846 19332
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16816 19264 16957 19292
rect 16816 19252 16822 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 18138 19292 18144 19304
rect 18099 19264 18144 19292
rect 16945 19255 17003 19261
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19292 18659 19295
rect 19150 19292 19156 19304
rect 18647 19264 19156 19292
rect 18647 19261 18659 19264
rect 18601 19255 18659 19261
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 17218 19224 17224 19236
rect 16684 19196 17224 19224
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 19720 19224 19748 19323
rect 19812 19292 19840 19323
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 19944 19332 19989 19360
rect 19944 19320 19950 19332
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20530 19360 20536 19372
rect 20128 19332 20173 19360
rect 20491 19332 20536 19360
rect 20128 19320 20134 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20626 19363 20684 19369
rect 20626 19329 20638 19363
rect 20672 19329 20684 19363
rect 20806 19360 20812 19372
rect 20767 19332 20812 19360
rect 20626 19323 20684 19329
rect 20254 19292 20260 19304
rect 19812 19264 20260 19292
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20548 19224 20576 19320
rect 19720 19196 20576 19224
rect 12066 19156 12072 19168
rect 12027 19128 12072 19156
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 12676 19128 13553 19156
rect 12676 19116 12682 19128
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 15562 19156 15568 19168
rect 15523 19128 15568 19156
rect 13541 19119 13599 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 16632 19128 17417 19156
rect 16632 19116 16638 19128
rect 17405 19125 17417 19128
rect 17451 19125 17463 19159
rect 17405 19119 17463 19125
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20640 19156 20668 19323
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 20990 19360 20996 19372
rect 20949 19332 20996 19360
rect 20990 19320 20996 19332
rect 21048 19369 21054 19372
rect 21048 19363 21097 19369
rect 21048 19329 21051 19363
rect 21085 19360 21097 19363
rect 21542 19360 21548 19372
rect 21085 19332 21548 19360
rect 21085 19329 21097 19332
rect 21048 19323 21097 19329
rect 21048 19320 21054 19323
rect 21542 19320 21548 19332
rect 21600 19320 21606 19372
rect 22830 19369 22836 19372
rect 22824 19360 22836 19369
rect 22791 19332 22836 19360
rect 22824 19323 22836 19332
rect 22830 19320 22836 19323
rect 22888 19320 22894 19372
rect 23566 19320 23572 19372
rect 23624 19360 23630 19372
rect 24673 19363 24731 19369
rect 24673 19360 24685 19363
rect 23624 19332 24685 19360
rect 23624 19320 23630 19332
rect 24673 19329 24685 19332
rect 24719 19360 24731 19363
rect 24762 19360 24768 19372
rect 24719 19332 24768 19360
rect 24719 19329 24731 19332
rect 24673 19323 24731 19329
rect 24762 19320 24768 19332
rect 24820 19320 24826 19372
rect 25406 19360 25412 19372
rect 25367 19332 25412 19360
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 22097 19295 22155 19301
rect 22097 19261 22109 19295
rect 22143 19292 22155 19295
rect 22554 19292 22560 19304
rect 22143 19264 22560 19292
rect 22143 19261 22155 19264
rect 22097 19255 22155 19261
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 25685 19295 25743 19301
rect 25685 19261 25697 19295
rect 25731 19292 25743 19295
rect 25866 19292 25872 19304
rect 25731 19264 25872 19292
rect 25731 19261 25743 19264
rect 25685 19255 25743 19261
rect 25866 19252 25872 19264
rect 25924 19252 25930 19304
rect 26206 19224 26234 19400
rect 27522 19360 27528 19372
rect 27483 19332 27528 19360
rect 27522 19320 27528 19332
rect 27580 19360 27586 19372
rect 28331 19363 28389 19369
rect 28331 19360 28343 19363
rect 27580 19332 28343 19360
rect 27580 19320 27586 19332
rect 28331 19329 28343 19332
rect 28377 19329 28389 19363
rect 28552 19335 28580 19400
rect 28810 19388 28816 19440
rect 28868 19428 28874 19440
rect 30193 19431 30251 19437
rect 30193 19428 30205 19431
rect 28868 19400 30205 19428
rect 28868 19388 28874 19400
rect 30193 19397 30205 19400
rect 30239 19397 30251 19431
rect 30193 19391 30251 19397
rect 30374 19388 30380 19440
rect 30432 19428 30438 19440
rect 30926 19428 30932 19440
rect 30432 19400 30932 19428
rect 30432 19388 30438 19400
rect 30926 19388 30932 19400
rect 30984 19388 30990 19440
rect 32858 19428 32864 19440
rect 32771 19400 32864 19428
rect 32858 19388 32864 19400
rect 32916 19428 32922 19440
rect 34790 19428 34796 19440
rect 32916 19400 34796 19428
rect 32916 19388 32922 19400
rect 34790 19388 34796 19400
rect 34848 19388 34854 19440
rect 29362 19360 29368 19372
rect 28331 19323 28389 19329
rect 28537 19329 28595 19335
rect 29323 19332 29368 19360
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19261 27215 19295
rect 27157 19255 27215 19261
rect 27249 19295 27307 19301
rect 27249 19261 27261 19295
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 27172 19224 27200 19255
rect 26206 19196 27200 19224
rect 20128 19128 20668 19156
rect 20128 19116 20134 19128
rect 23750 19116 23756 19168
rect 23808 19156 23814 19168
rect 23937 19159 23995 19165
rect 23937 19156 23949 19159
rect 23808 19128 23949 19156
rect 23808 19116 23814 19128
rect 23937 19125 23949 19128
rect 23983 19125 23995 19159
rect 23937 19119 23995 19125
rect 24026 19116 24032 19168
rect 24084 19156 24090 19168
rect 27264 19156 27292 19255
rect 27614 19252 27620 19304
rect 27672 19292 27678 19304
rect 28253 19295 28311 19301
rect 28253 19292 28265 19295
rect 27672 19264 28265 19292
rect 27672 19252 27678 19264
rect 28253 19261 28265 19264
rect 28299 19261 28311 19295
rect 28253 19255 28311 19261
rect 28445 19295 28503 19301
rect 28445 19261 28457 19295
rect 28491 19261 28503 19295
rect 28537 19295 28549 19329
rect 28583 19295 28595 19329
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 29546 19360 29552 19372
rect 29507 19332 29552 19360
rect 29546 19320 29552 19332
rect 29604 19320 29610 19372
rect 30834 19360 30840 19372
rect 30795 19332 30840 19360
rect 30834 19320 30840 19332
rect 30892 19320 30898 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 33689 19363 33747 19369
rect 33689 19360 33701 19363
rect 32456 19332 33701 19360
rect 32456 19320 32462 19332
rect 33689 19329 33701 19332
rect 33735 19329 33747 19363
rect 33689 19323 33747 19329
rect 28537 19289 28595 19295
rect 29638 19292 29644 19304
rect 29599 19264 29644 19292
rect 28445 19255 28503 19261
rect 28460 19156 28488 19255
rect 29638 19252 29644 19264
rect 29696 19252 29702 19304
rect 33134 19292 33140 19304
rect 33095 19264 33140 19292
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 28626 19184 28632 19236
rect 28684 19224 28690 19236
rect 30374 19224 30380 19236
rect 28684 19196 30380 19224
rect 28684 19184 28690 19196
rect 30374 19184 30380 19196
rect 30432 19184 30438 19236
rect 29178 19156 29184 19168
rect 24084 19128 28488 19156
rect 29139 19128 29184 19156
rect 24084 19116 24090 19128
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 29730 19116 29736 19168
rect 29788 19156 29794 19168
rect 30929 19159 30987 19165
rect 30929 19156 30941 19159
rect 29788 19128 30941 19156
rect 29788 19116 29794 19128
rect 30929 19125 30941 19128
rect 30975 19125 30987 19159
rect 30929 19119 30987 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 13446 18952 13452 18964
rect 13407 18924 13452 18952
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 16390 18952 16396 18964
rect 16351 18924 16396 18952
rect 16390 18912 16396 18924
rect 16448 18912 16454 18964
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20073 18955 20131 18961
rect 20073 18952 20085 18955
rect 19944 18924 20085 18952
rect 19944 18912 19950 18924
rect 20073 18921 20085 18924
rect 20119 18921 20131 18955
rect 20898 18952 20904 18964
rect 20073 18915 20131 18921
rect 20641 18924 20904 18952
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 20641 18884 20669 18924
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 21177 18955 21235 18961
rect 21177 18921 21189 18955
rect 21223 18952 21235 18955
rect 22094 18952 22100 18964
rect 21223 18924 22100 18952
rect 21223 18921 21235 18924
rect 21177 18915 21235 18921
rect 22094 18912 22100 18924
rect 22152 18912 22158 18964
rect 23290 18952 23296 18964
rect 23251 18924 23296 18952
rect 23290 18912 23296 18924
rect 23348 18912 23354 18964
rect 26234 18952 26240 18964
rect 23400 18924 26240 18952
rect 15528 18856 20669 18884
rect 15528 18844 15534 18856
rect 20714 18844 20720 18896
rect 20772 18884 20778 18896
rect 22281 18887 22339 18893
rect 22281 18884 22293 18887
rect 20772 18856 22293 18884
rect 20772 18844 20778 18856
rect 22281 18853 22293 18856
rect 22327 18853 22339 18887
rect 22281 18847 22339 18853
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18816 16911 18819
rect 16942 18816 16948 18828
rect 16899 18788 16948 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17368 18788 17785 18816
rect 17368 18776 17374 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 21082 18816 21088 18828
rect 17920 18788 17965 18816
rect 19444 18788 19656 18816
rect 17920 18776 17926 18788
rect 19444 18760 19472 18788
rect 11422 18748 11428 18760
rect 11335 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18748 11486 18760
rect 12802 18748 12808 18760
rect 11480 18720 12808 18748
rect 11480 18708 11486 18720
rect 12802 18708 12808 18720
rect 12860 18748 12866 18760
rect 13722 18748 13728 18760
rect 12860 18720 13728 18748
rect 12860 18708 12866 18720
rect 13722 18708 13728 18720
rect 13780 18748 13786 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13780 18720 14105 18748
rect 13780 18708 13786 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 16574 18748 16580 18760
rect 16535 18720 16580 18748
rect 14093 18711 14151 18717
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 11670 18683 11728 18689
rect 11670 18680 11682 18683
rect 11112 18652 11682 18680
rect 11112 18640 11118 18652
rect 11670 18649 11682 18652
rect 11716 18649 11728 18683
rect 13354 18680 13360 18692
rect 13315 18652 13360 18680
rect 11670 18643 11728 18649
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 13814 18640 13820 18692
rect 13872 18680 13878 18692
rect 14338 18683 14396 18689
rect 14338 18680 14350 18683
rect 13872 18652 14350 18680
rect 13872 18640 13878 18652
rect 14338 18649 14350 18652
rect 14384 18649 14396 18683
rect 14338 18643 14396 18649
rect 15930 18640 15936 18692
rect 15988 18680 15994 18692
rect 16776 18680 16804 18711
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17276 18720 17509 18748
rect 17276 18708 17282 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17678 18748 17684 18760
rect 17639 18720 17684 18748
rect 17497 18711 17555 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18748 18107 18751
rect 18598 18748 18604 18760
rect 18095 18720 18604 18748
rect 18095 18717 18107 18720
rect 18049 18711 18107 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19426 18748 19432 18760
rect 19387 18720 19432 18748
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19522 18751 19580 18757
rect 19522 18717 19534 18751
rect 19568 18717 19580 18751
rect 19522 18711 19580 18717
rect 18506 18680 18512 18692
rect 15988 18652 18512 18680
rect 15988 18640 15994 18652
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 19537 18680 19565 18711
rect 19392 18652 19565 18680
rect 19392 18640 19398 18652
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 11848 18584 12817 18612
rect 11848 18572 11854 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 15470 18612 15476 18624
rect 15431 18584 15476 18612
rect 12805 18575 12863 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 17678 18612 17684 18624
rect 16908 18584 17684 18612
rect 16908 18572 16914 18584
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 19426 18612 19432 18624
rect 18279 18584 19432 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 19628 18612 19656 18788
rect 19720 18788 21088 18816
rect 19720 18757 19748 18788
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 23400 18816 23428 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 27433 18955 27491 18961
rect 27433 18921 27445 18955
rect 27479 18952 27491 18955
rect 27614 18952 27620 18964
rect 27479 18924 27620 18952
rect 27479 18921 27491 18924
rect 27433 18915 27491 18921
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 29638 18912 29644 18964
rect 29696 18952 29702 18964
rect 30009 18955 30067 18961
rect 30009 18952 30021 18955
rect 29696 18924 30021 18952
rect 29696 18912 29702 18924
rect 30009 18921 30021 18924
rect 30055 18921 30067 18955
rect 30009 18915 30067 18921
rect 30282 18912 30288 18964
rect 30340 18952 30346 18964
rect 31113 18955 31171 18961
rect 31113 18952 31125 18955
rect 30340 18924 31125 18952
rect 30340 18912 30346 18924
rect 31113 18921 31125 18924
rect 31159 18921 31171 18955
rect 31113 18915 31171 18921
rect 32125 18955 32183 18961
rect 32125 18921 32137 18955
rect 32171 18952 32183 18955
rect 32214 18952 32220 18964
rect 32171 18924 32220 18952
rect 32171 18921 32183 18924
rect 32125 18915 32183 18921
rect 32214 18912 32220 18924
rect 32272 18912 32278 18964
rect 33318 18912 33324 18964
rect 33376 18952 33382 18964
rect 33873 18955 33931 18961
rect 33873 18952 33885 18955
rect 33376 18924 33885 18952
rect 33376 18912 33382 18924
rect 33873 18921 33885 18924
rect 33919 18921 33931 18955
rect 33873 18915 33931 18921
rect 23566 18884 23572 18896
rect 23527 18856 23572 18884
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 23658 18844 23664 18896
rect 23716 18884 23722 18896
rect 23716 18856 23761 18884
rect 23716 18844 23722 18856
rect 25222 18844 25228 18896
rect 25280 18884 25286 18896
rect 29454 18884 29460 18896
rect 25280 18856 25636 18884
rect 25280 18844 25286 18856
rect 24026 18816 24032 18828
rect 21600 18788 23428 18816
rect 23492 18788 24032 18816
rect 21600 18776 21606 18788
rect 19978 18757 19984 18760
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19935 18751 19984 18757
rect 19935 18717 19947 18751
rect 19981 18717 19984 18751
rect 19935 18711 19984 18717
rect 19978 18708 19984 18711
rect 20036 18708 20042 18760
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 19794 18680 19800 18692
rect 19755 18652 19800 18680
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 20548 18612 20576 18711
rect 20622 18708 20628 18760
rect 20680 18748 20686 18760
rect 20680 18720 20725 18748
rect 20680 18708 20686 18720
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20864 18720 20909 18748
rect 20864 18708 20870 18720
rect 20990 18708 20996 18760
rect 21048 18757 21054 18760
rect 21048 18748 21056 18757
rect 21634 18748 21640 18760
rect 21048 18720 21093 18748
rect 21595 18720 21640 18748
rect 21048 18711 21056 18720
rect 21048 18708 21054 18711
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 21744 18757 21772 18788
rect 21730 18751 21788 18757
rect 21730 18717 21742 18751
rect 21776 18717 21788 18751
rect 21730 18711 21788 18717
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 22143 18751 22201 18757
rect 22143 18717 22155 18751
rect 22189 18748 22201 18751
rect 22462 18748 22468 18760
rect 22189 18720 22468 18748
rect 22189 18717 22201 18720
rect 22143 18711 22201 18717
rect 20898 18680 20904 18692
rect 20859 18652 20904 18680
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 21928 18680 21956 18711
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 23492 18757 23520 18788
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 25314 18816 25320 18828
rect 25275 18788 25320 18816
rect 25314 18776 25320 18788
rect 25372 18776 25378 18828
rect 25608 18825 25636 18856
rect 27632 18856 29460 18884
rect 25593 18819 25651 18825
rect 25593 18785 25605 18819
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 27154 18776 27160 18828
rect 27212 18816 27218 18828
rect 27632 18825 27660 18856
rect 29454 18844 29460 18856
rect 29512 18844 29518 18896
rect 32766 18844 32772 18896
rect 32824 18884 32830 18896
rect 32824 18856 33088 18884
rect 32824 18844 32830 18856
rect 27617 18819 27675 18825
rect 27617 18816 27629 18819
rect 27212 18788 27629 18816
rect 27212 18776 27218 18788
rect 27617 18785 27629 18788
rect 27663 18785 27675 18819
rect 27617 18779 27675 18785
rect 27801 18819 27859 18825
rect 27801 18785 27813 18819
rect 27847 18816 27859 18819
rect 27982 18816 27988 18828
rect 27847 18788 27988 18816
rect 27847 18785 27859 18788
rect 27801 18779 27859 18785
rect 27982 18776 27988 18788
rect 28040 18816 28046 18828
rect 29086 18816 29092 18828
rect 28040 18788 29092 18816
rect 28040 18776 28046 18788
rect 29086 18776 29092 18788
rect 29144 18776 29150 18828
rect 32309 18819 32367 18825
rect 30208 18788 31064 18816
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18717 23535 18751
rect 23750 18748 23756 18760
rect 23711 18720 23756 18748
rect 23477 18711 23535 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 25332 18748 25360 18776
rect 30208 18760 30236 18788
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 24811 18720 25360 18748
rect 26620 18720 26985 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 21100 18652 21956 18680
rect 22002 18683 22060 18689
rect 19628 18584 20576 18612
rect 20806 18572 20812 18624
rect 20864 18612 20870 18624
rect 21100 18612 21128 18652
rect 22002 18649 22014 18683
rect 22048 18680 22060 18683
rect 22048 18652 22232 18680
rect 22048 18649 22060 18652
rect 22002 18643 22060 18649
rect 22204 18624 22232 18652
rect 22922 18640 22928 18692
rect 22980 18680 22986 18692
rect 23198 18680 23204 18692
rect 22980 18652 23204 18680
rect 22980 18640 22986 18652
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 24578 18680 24584 18692
rect 24539 18652 24584 18680
rect 24578 18640 24584 18652
rect 24636 18640 24642 18692
rect 25041 18683 25099 18689
rect 25041 18649 25053 18683
rect 25087 18680 25099 18683
rect 25866 18680 25872 18692
rect 25087 18652 25872 18680
rect 25087 18649 25099 18652
rect 25041 18643 25099 18649
rect 25866 18640 25872 18652
rect 25924 18640 25930 18692
rect 26620 18624 26648 18720
rect 26973 18717 26985 18720
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 27893 18751 27951 18757
rect 27764 18720 27809 18748
rect 27764 18708 27770 18720
rect 27893 18717 27905 18751
rect 27939 18748 27951 18751
rect 28074 18748 28080 18760
rect 27939 18720 28080 18748
rect 27939 18717 27951 18720
rect 27893 18711 27951 18717
rect 28074 18708 28080 18720
rect 28132 18708 28138 18760
rect 28350 18708 28356 18760
rect 28408 18748 28414 18760
rect 28445 18751 28503 18757
rect 28445 18748 28457 18751
rect 28408 18720 28457 18748
rect 28408 18708 28414 18720
rect 28445 18717 28457 18720
rect 28491 18717 28503 18751
rect 28718 18748 28724 18760
rect 28679 18720 28724 18748
rect 28445 18711 28503 18717
rect 28718 18708 28724 18720
rect 28776 18708 28782 18760
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18748 28871 18751
rect 29270 18748 29276 18760
rect 28859 18720 29276 18748
rect 28859 18717 28871 18720
rect 28813 18711 28871 18717
rect 29270 18708 29276 18720
rect 29328 18708 29334 18760
rect 30190 18748 30196 18760
rect 30151 18720 30196 18748
rect 30190 18708 30196 18720
rect 30248 18708 30254 18760
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18717 30343 18751
rect 30466 18748 30472 18760
rect 30427 18720 30472 18748
rect 30285 18711 30343 18717
rect 28166 18640 28172 18692
rect 28224 18680 28230 18692
rect 28629 18683 28687 18689
rect 28629 18680 28641 18683
rect 28224 18652 28641 18680
rect 28224 18640 28230 18652
rect 28629 18649 28641 18652
rect 28675 18649 28687 18683
rect 28629 18643 28687 18649
rect 30098 18640 30104 18692
rect 30156 18680 30162 18692
rect 30300 18680 30328 18711
rect 30466 18708 30472 18720
rect 30524 18708 30530 18760
rect 30558 18708 30564 18760
rect 30616 18748 30622 18760
rect 31036 18757 31064 18788
rect 32309 18785 32321 18819
rect 32355 18816 32367 18819
rect 33060 18816 33088 18856
rect 33226 18816 33232 18828
rect 32355 18788 32812 18816
rect 32355 18785 32367 18788
rect 32309 18779 32367 18785
rect 31021 18751 31079 18757
rect 30616 18720 30661 18748
rect 30616 18708 30622 18720
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31849 18751 31907 18757
rect 31849 18717 31861 18751
rect 31895 18748 31907 18751
rect 32030 18748 32036 18760
rect 31895 18720 32036 18748
rect 31895 18717 31907 18720
rect 31849 18711 31907 18717
rect 32030 18708 32036 18720
rect 32088 18708 32094 18760
rect 32784 18757 32812 18788
rect 33060 18788 33232 18816
rect 33060 18757 33088 18788
rect 33226 18776 33232 18788
rect 33284 18776 33290 18828
rect 32769 18751 32827 18757
rect 32769 18717 32781 18751
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18717 33103 18751
rect 33045 18711 33103 18717
rect 33134 18708 33140 18760
rect 33192 18748 33198 18760
rect 33781 18751 33839 18757
rect 33192 18720 33237 18748
rect 33192 18708 33198 18720
rect 33781 18717 33793 18751
rect 33827 18717 33839 18751
rect 33781 18711 33839 18717
rect 32950 18680 32956 18692
rect 30156 18652 30328 18680
rect 32911 18652 32956 18680
rect 30156 18640 30162 18652
rect 32950 18640 32956 18652
rect 33008 18640 33014 18692
rect 33796 18680 33824 18711
rect 33244 18652 33824 18680
rect 20864 18584 21128 18612
rect 20864 18572 20870 18584
rect 22186 18572 22192 18624
rect 22244 18572 22250 18624
rect 23106 18572 23112 18624
rect 23164 18612 23170 18624
rect 24854 18612 24860 18624
rect 23164 18584 24860 18612
rect 23164 18572 23170 18584
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 24949 18615 25007 18621
rect 24949 18581 24961 18615
rect 24995 18612 25007 18615
rect 25314 18612 25320 18624
rect 24995 18584 25320 18612
rect 24995 18581 25007 18584
rect 24949 18575 25007 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 26513 18615 26571 18621
rect 26513 18581 26525 18615
rect 26559 18612 26571 18615
rect 26602 18612 26608 18624
rect 26559 18584 26608 18612
rect 26559 18581 26571 18584
rect 26513 18575 26571 18581
rect 26602 18572 26608 18584
rect 26660 18572 26666 18624
rect 26789 18615 26847 18621
rect 26789 18581 26801 18615
rect 26835 18612 26847 18615
rect 27154 18612 27160 18624
rect 26835 18584 27160 18612
rect 26835 18581 26847 18584
rect 26789 18575 26847 18581
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 28994 18612 29000 18624
rect 28955 18584 29000 18612
rect 28994 18572 29000 18584
rect 29052 18572 29058 18624
rect 32582 18572 32588 18624
rect 32640 18612 32646 18624
rect 33244 18612 33272 18652
rect 32640 18584 33272 18612
rect 32640 18572 32646 18584
rect 33318 18572 33324 18624
rect 33376 18612 33382 18624
rect 33376 18584 33421 18612
rect 33376 18572 33382 18584
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 15010 18368 15016 18420
rect 15068 18408 15074 18420
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 15068 18380 15117 18408
rect 15068 18368 15074 18380
rect 15105 18377 15117 18380
rect 15151 18408 15163 18411
rect 15151 18380 19564 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 19536 18352 19564 18380
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 21266 18408 21272 18420
rect 20036 18380 21174 18408
rect 21227 18380 21272 18408
rect 20036 18368 20042 18380
rect 18138 18340 18144 18352
rect 15856 18312 18144 18340
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 11773 18275 11831 18281
rect 11773 18272 11785 18275
rect 10744 18244 11785 18272
rect 10744 18232 10750 18244
rect 11773 18241 11785 18244
rect 11819 18241 11831 18275
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 11773 18235 11831 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 13992 18275 14050 18281
rect 13992 18241 14004 18275
rect 14038 18272 14050 18275
rect 14550 18272 14556 18284
rect 14038 18244 14556 18272
rect 14038 18241 14050 18244
rect 13992 18235 14050 18241
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 15856 18281 15884 18312
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 19518 18300 19524 18352
rect 19576 18340 19582 18352
rect 20993 18343 21051 18349
rect 20993 18340 21005 18343
rect 19576 18312 21005 18340
rect 19576 18300 19582 18312
rect 20993 18309 21005 18312
rect 21039 18309 21051 18343
rect 20993 18303 21051 18309
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16025 18275 16083 18281
rect 16025 18272 16037 18275
rect 15988 18244 16037 18272
rect 15988 18232 15994 18244
rect 16025 18241 16037 18244
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 17957 18275 18015 18281
rect 17957 18272 17969 18275
rect 16264 18244 17969 18272
rect 16264 18232 16270 18244
rect 17957 18241 17969 18244
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 18224 18275 18282 18281
rect 18224 18241 18236 18275
rect 18270 18272 18282 18275
rect 19242 18272 19248 18284
rect 18270 18244 19248 18272
rect 18270 18241 18282 18244
rect 18224 18235 18282 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19628 18244 20177 18272
rect 11514 18204 11520 18216
rect 11475 18176 11520 18204
rect 11514 18164 11520 18176
rect 11572 18164 11578 18216
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18204 16911 18207
rect 16899 18176 16988 18204
rect 16899 18173 16911 18176
rect 16853 18167 16911 18173
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 12897 18071 12955 18077
rect 12897 18068 12909 18071
rect 12584 18040 12909 18068
rect 12584 18028 12590 18040
rect 12897 18037 12909 18040
rect 12943 18037 12955 18071
rect 12897 18031 12955 18037
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 15562 18068 15568 18080
rect 14516 18040 15568 18068
rect 14516 18028 14522 18040
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 15657 18071 15715 18077
rect 15657 18037 15669 18071
rect 15703 18068 15715 18071
rect 15746 18068 15752 18080
rect 15703 18040 15752 18068
rect 15703 18037 15715 18040
rect 15657 18031 15715 18037
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 16132 18068 16160 18167
rect 16960 18136 16988 18176
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 17092 18176 17141 18204
rect 17092 18164 17098 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 19058 18164 19064 18216
rect 19116 18204 19122 18216
rect 19628 18213 19656 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20718 18275 20776 18281
rect 20718 18241 20730 18275
rect 20764 18241 20776 18275
rect 20718 18235 20776 18241
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19116 18176 19625 18204
rect 19116 18164 19122 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 17954 18136 17960 18148
rect 16960 18108 17960 18136
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 20640 18136 20668 18235
rect 20733 18204 20761 18235
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21146 18281 21174 18380
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 22097 18411 22155 18417
rect 22097 18377 22109 18411
rect 22143 18408 22155 18411
rect 22278 18408 22284 18420
rect 22143 18380 22284 18408
rect 22143 18377 22155 18380
rect 22097 18371 22155 18377
rect 22278 18368 22284 18380
rect 22336 18368 22342 18420
rect 22462 18368 22468 18420
rect 22520 18368 22526 18420
rect 23014 18408 23020 18420
rect 22572 18380 23020 18408
rect 22480 18287 22508 18368
rect 21131 18275 21189 18281
rect 20956 18244 21001 18272
rect 20956 18232 20962 18244
rect 21131 18241 21143 18275
rect 21177 18272 21189 18275
rect 22002 18272 22008 18284
rect 21177 18244 22008 18272
rect 21177 18241 21189 18244
rect 21131 18235 21189 18241
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22462 18281 22520 18287
rect 22572 18281 22600 18380
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 25590 18408 25596 18420
rect 24320 18380 25596 18408
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18241 22431 18275
rect 22462 18247 22474 18281
rect 22508 18247 22520 18281
rect 22462 18241 22520 18247
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18241 22615 18275
rect 22373 18235 22431 18241
rect 22557 18235 22615 18241
rect 22741 18275 22799 18281
rect 22741 18241 22753 18275
rect 22787 18272 22799 18275
rect 22922 18272 22928 18284
rect 22787 18244 22928 18272
rect 22787 18241 22799 18244
rect 22741 18235 22799 18241
rect 21266 18204 21272 18216
rect 20733 18176 21272 18204
rect 20714 18136 20720 18148
rect 18892 18108 20576 18136
rect 20640 18108 20720 18136
rect 17034 18068 17040 18080
rect 16132 18040 17040 18068
rect 17034 18028 17040 18040
rect 17092 18068 17098 18080
rect 18892 18068 18920 18108
rect 17092 18040 18920 18068
rect 19337 18071 19395 18077
rect 17092 18028 17098 18040
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19518 18068 19524 18080
rect 19383 18040 19524 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19668 18040 19993 18068
rect 19668 18028 19674 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 20548 18068 20576 18108
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 20824 18068 20852 18176
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 22388 18204 22416 18235
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 24320 18281 24348 18380
rect 25590 18368 25596 18380
rect 25648 18408 25654 18420
rect 27341 18411 27399 18417
rect 27341 18408 27353 18411
rect 25648 18380 27353 18408
rect 25648 18368 25654 18380
rect 27341 18377 27353 18380
rect 27387 18408 27399 18411
rect 28074 18408 28080 18420
rect 27387 18380 28080 18408
rect 27387 18377 27399 18380
rect 27341 18371 27399 18377
rect 28074 18368 28080 18380
rect 28132 18368 28138 18420
rect 29181 18411 29239 18417
rect 29181 18377 29193 18411
rect 29227 18408 29239 18411
rect 29362 18408 29368 18420
rect 29227 18380 29368 18408
rect 29227 18377 29239 18380
rect 29181 18371 29239 18377
rect 29362 18368 29368 18380
rect 29420 18368 29426 18420
rect 30377 18411 30435 18417
rect 30377 18377 30389 18411
rect 30423 18408 30435 18411
rect 30558 18408 30564 18420
rect 30423 18380 30564 18408
rect 30423 18377 30435 18380
rect 30377 18371 30435 18377
rect 30558 18368 30564 18380
rect 30616 18368 30622 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 32490 18408 32496 18420
rect 30708 18380 32496 18408
rect 30708 18368 30714 18380
rect 32490 18368 32496 18380
rect 32548 18408 32554 18420
rect 33594 18408 33600 18420
rect 32548 18380 33600 18408
rect 32548 18368 32554 18380
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 25133 18343 25191 18349
rect 25133 18309 25145 18343
rect 25179 18340 25191 18343
rect 25222 18340 25228 18352
rect 25179 18312 25228 18340
rect 25179 18309 25191 18312
rect 25133 18303 25191 18309
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 26421 18343 26479 18349
rect 26421 18309 26433 18343
rect 26467 18340 26479 18343
rect 28258 18340 28264 18352
rect 26467 18312 28264 18340
rect 26467 18309 26479 18312
rect 26421 18303 26479 18309
rect 28258 18300 28264 18312
rect 28316 18300 28322 18352
rect 31018 18340 31024 18352
rect 30979 18312 31024 18340
rect 31018 18300 31024 18312
rect 31076 18300 31082 18352
rect 32398 18300 32404 18352
rect 32456 18340 32462 18352
rect 33686 18340 33692 18352
rect 32456 18312 33692 18340
rect 32456 18300 32462 18312
rect 33686 18300 33692 18312
rect 33744 18300 33750 18352
rect 33870 18300 33876 18352
rect 33928 18340 33934 18352
rect 33965 18343 34023 18349
rect 33965 18340 33977 18343
rect 33928 18312 33977 18340
rect 33928 18300 33934 18312
rect 33965 18309 33977 18312
rect 34011 18309 34023 18343
rect 33965 18303 34023 18309
rect 34154 18284 34212 18287
rect 23569 18275 23627 18281
rect 23569 18272 23581 18275
rect 23078 18244 23581 18272
rect 23078 18216 23106 18244
rect 23569 18241 23581 18244
rect 23615 18241 23627 18275
rect 23569 18235 23627 18241
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 22646 18204 22652 18216
rect 22388 18176 22652 18204
rect 22646 18164 22652 18176
rect 22704 18204 22710 18216
rect 22830 18204 22836 18216
rect 22704 18176 22836 18204
rect 22704 18164 22710 18176
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 23014 18164 23020 18216
rect 23072 18176 23106 18216
rect 23072 18164 23078 18176
rect 23198 18164 23204 18216
rect 23256 18204 23262 18216
rect 24412 18204 24440 18235
rect 24486 18232 24492 18284
rect 24544 18272 24550 18284
rect 24544 18244 24589 18272
rect 24544 18232 24550 18244
rect 24670 18232 24676 18284
rect 24728 18272 24734 18284
rect 25314 18272 25320 18284
rect 24728 18244 24773 18272
rect 25275 18244 25320 18272
rect 24728 18232 24734 18244
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18272 25467 18275
rect 25866 18272 25872 18284
rect 25455 18244 25872 18272
rect 25455 18241 25467 18244
rect 25409 18235 25467 18241
rect 25866 18232 25872 18244
rect 25924 18232 25930 18284
rect 26237 18275 26295 18281
rect 26237 18241 26249 18275
rect 26283 18241 26295 18275
rect 26237 18235 26295 18241
rect 23256 18176 24440 18204
rect 23256 18164 23262 18176
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 24578 18136 24584 18148
rect 20956 18108 24584 18136
rect 20956 18096 20962 18108
rect 24578 18096 24584 18108
rect 24636 18096 24642 18148
rect 24854 18096 24860 18148
rect 24912 18136 24918 18148
rect 25133 18139 25191 18145
rect 25133 18136 25145 18139
rect 24912 18108 25145 18136
rect 24912 18096 24918 18108
rect 25133 18105 25145 18108
rect 25179 18136 25191 18139
rect 25498 18136 25504 18148
rect 25179 18108 25504 18136
rect 25179 18105 25191 18108
rect 25133 18099 25191 18105
rect 25498 18096 25504 18108
rect 25556 18096 25562 18148
rect 26252 18136 26280 18235
rect 27062 18232 27068 18284
rect 27120 18272 27126 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 27120 18244 27169 18272
rect 27120 18232 27126 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18272 27307 18275
rect 27798 18272 27804 18284
rect 27295 18244 27804 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 27798 18232 27804 18244
rect 27856 18232 27862 18284
rect 27982 18272 27988 18284
rect 27943 18244 27988 18272
rect 27982 18232 27988 18244
rect 28040 18232 28046 18284
rect 28166 18272 28172 18284
rect 28127 18244 28172 18272
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18272 28595 18275
rect 28718 18272 28724 18284
rect 28583 18244 28724 18272
rect 28583 18241 28595 18244
rect 28537 18235 28595 18241
rect 28718 18232 28724 18244
rect 28776 18232 28782 18284
rect 29086 18232 29092 18284
rect 29144 18272 29150 18284
rect 29549 18275 29607 18281
rect 29549 18272 29561 18275
rect 29144 18244 29561 18272
rect 29144 18232 29150 18244
rect 29549 18241 29561 18244
rect 29595 18241 29607 18275
rect 29730 18272 29736 18284
rect 29691 18244 29736 18272
rect 29549 18235 29607 18241
rect 29730 18232 29736 18244
rect 29788 18232 29794 18284
rect 29917 18275 29975 18281
rect 29917 18241 29929 18275
rect 29963 18241 29975 18275
rect 29917 18235 29975 18241
rect 27525 18207 27583 18213
rect 27525 18173 27537 18207
rect 27571 18204 27583 18207
rect 28000 18204 28028 18232
rect 28258 18204 28264 18216
rect 27571 18176 28028 18204
rect 28219 18176 28264 18204
rect 27571 18173 27583 18176
rect 27525 18167 27583 18173
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18204 28411 18207
rect 29270 18204 29276 18216
rect 28399 18176 29276 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 29270 18164 29276 18176
rect 29328 18164 29334 18216
rect 29932 18204 29960 18235
rect 30282 18232 30288 18284
rect 30340 18272 30346 18284
rect 30653 18275 30711 18281
rect 30653 18272 30665 18275
rect 30340 18244 30665 18272
rect 30340 18232 30346 18244
rect 30653 18241 30665 18244
rect 30699 18241 30711 18275
rect 30926 18272 30932 18284
rect 30887 18244 30932 18272
rect 30653 18235 30711 18241
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 32582 18232 32588 18284
rect 32640 18272 32646 18284
rect 32953 18275 33011 18281
rect 32953 18272 32965 18275
rect 32640 18244 32965 18272
rect 32640 18232 32646 18244
rect 32953 18241 32965 18244
rect 32999 18241 33011 18275
rect 32953 18235 33011 18241
rect 33045 18275 33103 18281
rect 33045 18241 33057 18275
rect 33091 18241 33103 18275
rect 33045 18235 33103 18241
rect 30098 18204 30104 18216
rect 29932 18176 30104 18204
rect 30098 18164 30104 18176
rect 30156 18204 30162 18216
rect 30561 18207 30619 18213
rect 30561 18204 30573 18207
rect 30156 18176 30573 18204
rect 30156 18164 30162 18176
rect 30561 18173 30573 18176
rect 30607 18173 30619 18207
rect 30561 18167 30619 18173
rect 32858 18164 32864 18216
rect 32916 18204 32922 18216
rect 33060 18204 33088 18235
rect 33226 18232 33232 18284
rect 33284 18272 33290 18284
rect 33321 18275 33379 18281
rect 33321 18272 33333 18275
rect 33284 18244 33333 18272
rect 33284 18232 33290 18244
rect 33321 18241 33333 18244
rect 33367 18241 33379 18275
rect 33321 18235 33379 18241
rect 32916 18176 33088 18204
rect 33336 18204 33364 18235
rect 33594 18232 33600 18284
rect 33652 18272 33658 18284
rect 33781 18275 33839 18281
rect 33781 18272 33793 18275
rect 33652 18244 33793 18272
rect 33652 18232 33658 18244
rect 33781 18241 33793 18244
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 34057 18275 34115 18281
rect 34057 18241 34069 18275
rect 34103 18241 34115 18275
rect 34057 18235 34115 18241
rect 34072 18204 34100 18235
rect 34146 18232 34152 18284
rect 34204 18278 34212 18284
rect 34204 18250 34243 18278
rect 34204 18241 34212 18250
rect 34204 18232 34210 18241
rect 33336 18176 34100 18204
rect 32916 18164 32922 18176
rect 27614 18136 27620 18148
rect 26252 18108 27620 18136
rect 27614 18096 27620 18108
rect 27672 18096 27678 18148
rect 28902 18096 28908 18148
rect 28960 18136 28966 18148
rect 29457 18139 29515 18145
rect 29457 18136 29469 18139
rect 28960 18108 29469 18136
rect 28960 18096 28966 18108
rect 29457 18105 29469 18108
rect 29503 18105 29515 18139
rect 29457 18099 29515 18105
rect 29641 18139 29699 18145
rect 29641 18105 29653 18139
rect 29687 18136 29699 18139
rect 30926 18136 30932 18148
rect 29687 18108 30932 18136
rect 29687 18105 29699 18108
rect 29641 18099 29699 18105
rect 30926 18096 30932 18108
rect 30984 18096 30990 18148
rect 31386 18096 31392 18148
rect 31444 18136 31450 18148
rect 33781 18139 33839 18145
rect 33781 18136 33793 18139
rect 31444 18108 33793 18136
rect 31444 18096 31450 18108
rect 33781 18105 33793 18108
rect 33827 18105 33839 18139
rect 33781 18099 33839 18105
rect 20548 18040 20852 18068
rect 19981 18031 20039 18037
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 23014 18068 23020 18080
rect 22428 18040 23020 18068
rect 22428 18028 22434 18040
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 23382 18068 23388 18080
rect 23343 18040 23388 18068
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 24029 18071 24087 18077
rect 24029 18037 24041 18071
rect 24075 18068 24087 18071
rect 24946 18068 24952 18080
rect 24075 18040 24952 18068
rect 24075 18037 24087 18040
rect 24029 18031 24087 18037
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18068 27491 18071
rect 27522 18068 27528 18080
rect 27479 18040 27528 18068
rect 27479 18037 27491 18040
rect 27433 18031 27491 18037
rect 27522 18028 27528 18040
rect 27580 18028 27586 18080
rect 28721 18071 28779 18077
rect 28721 18037 28733 18071
rect 28767 18068 28779 18071
rect 29362 18068 29368 18080
rect 28767 18040 29368 18068
rect 28767 18037 28779 18040
rect 28721 18031 28779 18037
rect 29362 18028 29368 18040
rect 29420 18028 29426 18080
rect 31754 18028 31760 18080
rect 31812 18068 31818 18080
rect 32769 18071 32827 18077
rect 32769 18068 32781 18071
rect 31812 18040 32781 18068
rect 31812 18028 31818 18040
rect 32769 18037 32781 18040
rect 32815 18068 32827 18071
rect 32950 18068 32956 18080
rect 32815 18040 32956 18068
rect 32815 18037 32827 18040
rect 32769 18031 32827 18037
rect 32950 18028 32956 18040
rect 33008 18028 33014 18080
rect 33134 18028 33140 18080
rect 33192 18068 33198 18080
rect 33229 18071 33287 18077
rect 33229 18068 33241 18071
rect 33192 18040 33241 18068
rect 33192 18028 33198 18040
rect 33229 18037 33241 18040
rect 33275 18068 33287 18071
rect 34146 18068 34152 18080
rect 33275 18040 34152 18068
rect 33275 18037 33287 18040
rect 33229 18031 33287 18037
rect 34146 18028 34152 18040
rect 34204 18028 34210 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11790 17864 11796 17876
rect 10827 17836 11796 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 14550 17864 14556 17876
rect 14511 17836 14556 17864
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 16850 17864 16856 17876
rect 14752 17836 16856 17864
rect 14752 17796 14780 17836
rect 16850 17824 16856 17836
rect 16908 17824 16914 17876
rect 17034 17864 17040 17876
rect 16995 17836 17040 17864
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 18196 17836 18245 17864
rect 18196 17824 18202 17836
rect 18233 17833 18245 17836
rect 18279 17833 18291 17867
rect 19242 17864 19248 17876
rect 19203 17836 19248 17864
rect 18233 17827 18291 17833
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 21174 17864 21180 17876
rect 21135 17836 21180 17864
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 22189 17867 22247 17873
rect 22189 17833 22201 17867
rect 22235 17833 22247 17867
rect 22189 17827 22247 17833
rect 13556 17768 14780 17796
rect 11422 17728 11428 17740
rect 11383 17700 11428 17728
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 13556 17737 13584 17768
rect 18506 17756 18512 17808
rect 18564 17796 18570 17808
rect 19613 17799 19671 17805
rect 19613 17796 19625 17799
rect 18564 17768 19625 17796
rect 18564 17756 18570 17768
rect 19613 17765 19625 17768
rect 19659 17765 19671 17799
rect 19613 17759 19671 17765
rect 20806 17756 20812 17808
rect 20864 17756 20870 17808
rect 22204 17796 22232 17827
rect 28074 17824 28080 17876
rect 28132 17864 28138 17876
rect 28169 17867 28227 17873
rect 28169 17864 28181 17867
rect 28132 17836 28181 17864
rect 28132 17824 28138 17836
rect 28169 17833 28181 17836
rect 28215 17833 28227 17867
rect 28169 17827 28227 17833
rect 28813 17867 28871 17873
rect 28813 17833 28825 17867
rect 28859 17864 28871 17867
rect 29178 17864 29184 17876
rect 28859 17836 29184 17864
rect 28859 17833 28871 17836
rect 28813 17827 28871 17833
rect 29178 17824 29184 17836
rect 29236 17824 29242 17876
rect 29638 17824 29644 17876
rect 29696 17864 29702 17876
rect 29917 17867 29975 17873
rect 29917 17864 29929 17867
rect 29696 17836 29929 17864
rect 29696 17824 29702 17836
rect 29917 17833 29929 17836
rect 29963 17833 29975 17867
rect 33318 17864 33324 17876
rect 29917 17827 29975 17833
rect 30392 17836 33324 17864
rect 23106 17796 23112 17808
rect 22204 17768 23112 17796
rect 23106 17756 23112 17768
rect 23164 17756 23170 17808
rect 27798 17756 27804 17808
rect 27856 17796 27862 17808
rect 28905 17799 28963 17805
rect 28905 17796 28917 17799
rect 27856 17768 28917 17796
rect 27856 17756 27862 17768
rect 28905 17765 28917 17768
rect 28951 17765 28963 17799
rect 30392 17796 30420 17836
rect 33318 17824 33324 17836
rect 33376 17824 33382 17876
rect 28905 17759 28963 17765
rect 29012 17768 30420 17796
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17697 13599 17731
rect 15010 17728 15016 17740
rect 14971 17700 15016 17728
rect 13541 17691 13599 17697
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 17862 17728 17868 17740
rect 17823 17700 17868 17728
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 19518 17688 19524 17740
rect 19576 17728 19582 17740
rect 19576 17700 19748 17728
rect 19576 17688 19582 17700
rect 11692 17663 11750 17669
rect 11692 17629 11704 17663
rect 11738 17660 11750 17663
rect 12066 17660 12072 17672
rect 11738 17632 12072 17660
rect 11738 17629 11750 17632
rect 11692 17623 11750 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 14550 17660 14556 17672
rect 13403 17632 14556 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17660 14979 17663
rect 15102 17660 15108 17672
rect 14967 17632 15108 17660
rect 14967 17629 14979 17632
rect 14921 17623 14979 17629
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 15657 17663 15715 17669
rect 15657 17629 15669 17663
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 10594 17592 10600 17604
rect 10555 17564 10600 17592
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 10813 17595 10871 17601
rect 10813 17561 10825 17595
rect 10859 17592 10871 17595
rect 11606 17592 11612 17604
rect 10859 17564 11612 17592
rect 10859 17561 10871 17564
rect 10813 17555 10871 17561
rect 11606 17552 11612 17564
rect 11664 17552 11670 17604
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 15378 17592 15384 17604
rect 13780 17564 15384 17592
rect 13780 17552 13786 17564
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 15672 17592 15700 17623
rect 15746 17620 15752 17672
rect 15804 17660 15810 17672
rect 15924 17663 15982 17669
rect 15924 17660 15936 17663
rect 15804 17632 15936 17660
rect 15804 17620 15810 17632
rect 15924 17629 15936 17632
rect 15970 17629 15982 17663
rect 15924 17623 15982 17629
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17497 17663 17555 17669
rect 17497 17660 17509 17663
rect 17276 17632 17509 17660
rect 17276 17620 17282 17632
rect 17497 17629 17509 17632
rect 17543 17629 17555 17663
rect 17678 17660 17684 17672
rect 17639 17632 17684 17660
rect 17497 17623 17555 17629
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 18049 17663 18107 17669
rect 18049 17629 18061 17663
rect 18095 17660 18107 17663
rect 18874 17660 18880 17672
rect 18095 17632 18880 17660
rect 18095 17629 18107 17632
rect 18049 17623 18107 17629
rect 16206 17592 16212 17604
rect 15672 17564 16212 17592
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 10962 17524 10968 17536
rect 10923 17496 10968 17524
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 11756 17496 12817 17524
rect 11756 17484 11762 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 12805 17487 12863 17493
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 17218 17524 17224 17536
rect 14608 17496 17224 17524
rect 14608 17484 14614 17496
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17788 17524 17816 17623
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19720 17669 19748 17700
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20070 17660 20076 17672
rect 19751 17632 20076 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20530 17660 20536 17672
rect 20491 17632 20536 17660
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 20626 17663 20684 17669
rect 20626 17629 20638 17663
rect 20672 17660 20684 17663
rect 20714 17660 20720 17672
rect 20672 17632 20720 17660
rect 20672 17629 20684 17632
rect 20626 17623 20684 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 20824 17669 20852 17756
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 23198 17728 23204 17740
rect 22520 17700 23204 17728
rect 22520 17688 22526 17700
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 20990 17620 20996 17672
rect 21048 17669 21054 17672
rect 21048 17660 21056 17669
rect 22922 17660 22928 17672
rect 21048 17632 21093 17660
rect 22883 17632 22928 17660
rect 21048 17623 21056 17632
rect 21048 17620 21054 17623
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 23032 17669 23060 17700
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 26786 17728 26792 17740
rect 26747 17700 26792 17728
rect 26786 17688 26792 17700
rect 26844 17688 26850 17740
rect 29012 17737 29040 17768
rect 30466 17756 30472 17808
rect 30524 17796 30530 17808
rect 30653 17799 30711 17805
rect 30653 17796 30665 17799
rect 30524 17768 30665 17796
rect 30524 17756 30530 17768
rect 30653 17765 30665 17768
rect 30699 17765 30711 17799
rect 30653 17759 30711 17765
rect 31481 17799 31539 17805
rect 31481 17765 31493 17799
rect 31527 17765 31539 17799
rect 32030 17796 32036 17808
rect 31943 17768 32036 17796
rect 31481 17759 31539 17765
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17697 29055 17731
rect 31496 17728 31524 17759
rect 32030 17756 32036 17768
rect 32088 17796 32094 17808
rect 33229 17799 33287 17805
rect 33229 17796 33241 17799
rect 32088 17768 33241 17796
rect 32088 17756 32094 17768
rect 33229 17765 33241 17768
rect 33275 17765 33287 17799
rect 33229 17759 33287 17765
rect 31754 17728 31760 17740
rect 28997 17691 29055 17697
rect 29288 17700 31524 17728
rect 31715 17700 31760 17728
rect 23017 17663 23075 17669
rect 23017 17629 23029 17663
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 23164 17632 23209 17660
rect 23164 17620 23170 17632
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23566 17660 23572 17672
rect 23348 17632 23572 17660
rect 23348 17620 23354 17632
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 24854 17660 24860 17672
rect 24815 17632 24860 17660
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 24946 17620 24952 17672
rect 25004 17660 25010 17672
rect 27045 17663 27103 17669
rect 27045 17660 27057 17663
rect 25004 17632 27057 17660
rect 25004 17620 25010 17632
rect 27045 17629 27057 17632
rect 27091 17629 27103 17663
rect 27045 17623 27103 17629
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17660 28779 17663
rect 29288 17660 29316 17700
rect 28767 17632 29316 17660
rect 28767 17629 28779 17632
rect 28721 17623 28779 17629
rect 29362 17620 29368 17672
rect 29420 17660 29426 17672
rect 29932 17669 29960 17700
rect 31754 17688 31760 17700
rect 31812 17688 31818 17740
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 29420 17632 29561 17660
rect 29420 17620 29426 17632
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 29917 17663 29975 17669
rect 29917 17629 29929 17663
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 30101 17663 30159 17669
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 30653 17663 30711 17669
rect 30653 17629 30665 17663
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 30837 17663 30895 17669
rect 30837 17629 30849 17663
rect 30883 17660 30895 17663
rect 30926 17660 30932 17672
rect 30883 17632 30932 17660
rect 30883 17629 30895 17632
rect 30837 17623 30895 17629
rect 20901 17595 20959 17601
rect 20901 17561 20913 17595
rect 20947 17592 20959 17595
rect 21174 17592 21180 17604
rect 20947 17564 21180 17592
rect 20947 17561 20959 17564
rect 20901 17555 20959 17561
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 21821 17595 21879 17601
rect 21821 17592 21833 17595
rect 21692 17564 21833 17592
rect 21692 17552 21698 17564
rect 21821 17561 21833 17564
rect 21867 17561 21879 17595
rect 21821 17555 21879 17561
rect 22005 17595 22063 17601
rect 22005 17561 22017 17595
rect 22051 17561 22063 17595
rect 22005 17555 22063 17561
rect 17552 17496 17816 17524
rect 17552 17484 17558 17496
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 22020 17524 22048 17555
rect 24578 17552 24584 17604
rect 24636 17592 24642 17604
rect 25102 17595 25160 17601
rect 25102 17592 25114 17595
rect 24636 17564 25114 17592
rect 24636 17552 24642 17564
rect 25102 17561 25114 17564
rect 25148 17561 25160 17595
rect 25102 17555 25160 17561
rect 25590 17552 25596 17604
rect 25648 17592 25654 17604
rect 26050 17592 26056 17604
rect 25648 17564 26056 17592
rect 25648 17552 25654 17564
rect 26050 17552 26056 17564
rect 26108 17552 26114 17604
rect 29086 17552 29092 17604
rect 29144 17592 29150 17604
rect 30116 17592 30144 17623
rect 29144 17564 30144 17592
rect 30668 17592 30696 17623
rect 30926 17620 30932 17632
rect 30984 17620 30990 17672
rect 31386 17660 31392 17672
rect 31347 17632 31392 17660
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 31018 17592 31024 17604
rect 30668 17564 31024 17592
rect 29144 17552 29150 17564
rect 31018 17552 31024 17564
rect 31076 17552 31082 17604
rect 31481 17595 31539 17601
rect 31481 17561 31493 17595
rect 31527 17592 31539 17595
rect 32048 17592 32076 17756
rect 32214 17728 32220 17740
rect 32175 17700 32220 17728
rect 32214 17688 32220 17700
rect 32272 17688 32278 17740
rect 32677 17731 32735 17737
rect 32677 17697 32689 17731
rect 32723 17728 32735 17731
rect 33410 17728 33416 17740
rect 32723 17700 33416 17728
rect 32723 17697 32735 17700
rect 32677 17691 32735 17697
rect 33410 17688 33416 17700
rect 33468 17688 33474 17740
rect 32398 17660 32404 17672
rect 32359 17632 32404 17660
rect 32398 17620 32404 17632
rect 32456 17620 32462 17672
rect 32490 17620 32496 17672
rect 32548 17660 32554 17672
rect 32766 17660 32772 17672
rect 32548 17632 32593 17660
rect 32727 17632 32772 17660
rect 32548 17620 32554 17632
rect 32766 17620 32772 17632
rect 32824 17660 32830 17672
rect 32824 17632 33180 17660
rect 32824 17620 32830 17632
rect 31527 17564 32076 17592
rect 33152 17592 33180 17632
rect 33594 17620 33600 17672
rect 33652 17669 33658 17672
rect 33652 17660 33660 17669
rect 33652 17632 33697 17660
rect 33652 17623 33660 17632
rect 33652 17620 33658 17623
rect 33229 17595 33287 17601
rect 33229 17592 33241 17595
rect 33152 17564 33241 17592
rect 31527 17561 31539 17564
rect 31481 17555 31539 17561
rect 33229 17561 33241 17564
rect 33275 17561 33287 17595
rect 33410 17592 33416 17604
rect 33371 17564 33416 17592
rect 33229 17555 33287 17561
rect 33410 17552 33416 17564
rect 33468 17552 33474 17604
rect 33505 17595 33563 17601
rect 33505 17561 33517 17595
rect 33551 17561 33563 17595
rect 33505 17555 33563 17561
rect 22646 17524 22652 17536
rect 21140 17496 22048 17524
rect 22607 17496 22652 17524
rect 21140 17484 21146 17496
rect 22646 17484 22652 17496
rect 22704 17484 22710 17536
rect 24762 17484 24768 17536
rect 24820 17524 24826 17536
rect 25866 17524 25872 17536
rect 24820 17496 25872 17524
rect 24820 17484 24826 17496
rect 25866 17484 25872 17496
rect 25924 17524 25930 17536
rect 26237 17527 26295 17533
rect 26237 17524 26249 17527
rect 25924 17496 26249 17524
rect 25924 17484 25930 17496
rect 26237 17493 26249 17496
rect 26283 17493 26295 17527
rect 26237 17487 26295 17493
rect 29454 17484 29460 17536
rect 29512 17524 29518 17536
rect 29733 17527 29791 17533
rect 29733 17524 29745 17527
rect 29512 17496 29745 17524
rect 29512 17484 29518 17496
rect 29733 17493 29745 17496
rect 29779 17493 29791 17527
rect 29733 17487 29791 17493
rect 31573 17527 31631 17533
rect 31573 17493 31585 17527
rect 31619 17524 31631 17527
rect 32214 17524 32220 17536
rect 31619 17496 32220 17524
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 32214 17484 32220 17496
rect 32272 17484 32278 17536
rect 32858 17484 32864 17536
rect 32916 17524 32922 17536
rect 33520 17524 33548 17555
rect 32916 17496 33548 17524
rect 32916 17484 32922 17496
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12555 17323 12613 17329
rect 12555 17320 12567 17323
rect 11940 17292 11985 17320
rect 12268 17292 12567 17320
rect 11940 17280 11946 17292
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 11517 17255 11575 17261
rect 11517 17252 11529 17255
rect 10652 17224 11529 17252
rect 10652 17212 10658 17224
rect 11517 17221 11529 17224
rect 11563 17221 11575 17255
rect 11517 17215 11575 17221
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11532 17184 11560 17215
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 11733 17255 11791 17261
rect 11733 17252 11745 17255
rect 11664 17224 11745 17252
rect 11664 17212 11670 17224
rect 11733 17221 11745 17224
rect 11779 17252 11791 17255
rect 12268 17252 12296 17292
rect 12555 17289 12567 17292
rect 12601 17320 12613 17323
rect 12986 17320 12992 17332
rect 12601 17292 12992 17320
rect 12601 17289 12613 17292
rect 12555 17283 12613 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13633 17323 13691 17329
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13814 17320 13820 17332
rect 13679 17292 13820 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14458 17320 14464 17332
rect 13924 17292 14464 17320
rect 11779 17224 12296 17252
rect 12391 17255 12449 17261
rect 11779 17221 11791 17224
rect 11733 17215 11791 17221
rect 12391 17221 12403 17255
rect 12437 17252 12449 17255
rect 12894 17252 12900 17264
rect 12437 17224 12900 17252
rect 12437 17221 12449 17224
rect 12391 17215 12449 17221
rect 12406 17184 12434 17215
rect 12894 17212 12900 17224
rect 12952 17252 12958 17264
rect 13924 17252 13952 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 14792 17292 15301 17320
rect 14792 17280 14798 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 24578 17320 24584 17332
rect 16163 17292 23106 17320
rect 24539 17292 24584 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 12952 17224 13952 17252
rect 12952 17212 12958 17224
rect 14366 17212 14372 17264
rect 14424 17252 14430 17264
rect 14424 17224 14780 17252
rect 14424 17212 14430 17224
rect 13814 17184 13820 17196
rect 11532 17156 12434 17184
rect 13775 17156 13820 17184
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14550 17184 14556 17196
rect 14056 17156 14556 17184
rect 14056 17144 14062 17156
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 14752 17193 14780 17224
rect 14826 17212 14832 17264
rect 14884 17252 14890 17264
rect 16761 17255 16819 17261
rect 14884 17224 15700 17252
rect 14884 17212 14890 17224
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 15068 17156 15117 17184
rect 15068 17144 15074 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 14093 17119 14151 17125
rect 14093 17085 14105 17119
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 10781 17051 10839 17057
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 11054 17048 11060 17060
rect 10827 17020 11060 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 12713 17051 12771 17057
rect 12713 17048 12725 17051
rect 11296 17020 12725 17048
rect 11296 17008 11302 17020
rect 12713 17017 12725 17020
rect 12759 17017 12771 17051
rect 14108 17048 14136 17079
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14700 17088 14841 17116
rect 14700 17076 14706 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 14918 17076 14924 17128
rect 14976 17116 14982 17128
rect 15672 17116 15700 17224
rect 16761 17221 16773 17255
rect 16807 17252 16819 17255
rect 17926 17255 17984 17261
rect 17926 17252 17938 17255
rect 16807 17224 17938 17252
rect 16807 17221 16819 17224
rect 16761 17215 16819 17221
rect 17926 17221 17938 17224
rect 17972 17221 17984 17255
rect 17926 17215 17984 17221
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 20622 17252 20628 17264
rect 19484 17224 20628 17252
rect 19484 17212 19490 17224
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 21266 17212 21272 17264
rect 21324 17252 21330 17264
rect 22186 17252 22192 17264
rect 21324 17224 22192 17252
rect 21324 17212 21330 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22646 17212 22652 17264
rect 22704 17252 22710 17264
rect 22986 17255 23044 17261
rect 22986 17252 22998 17255
rect 22704 17224 22998 17252
rect 22704 17212 22710 17224
rect 22986 17221 22998 17224
rect 23032 17221 23044 17255
rect 22986 17215 23044 17221
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 15933 17187 15991 17193
rect 15804 17156 15849 17184
rect 15804 17144 15810 17156
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 16022 17184 16028 17196
rect 15979 17156 16028 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 16942 17184 16948 17196
rect 16903 17156 16948 17184
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17126 17184 17132 17196
rect 17087 17156 17132 17184
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 19518 17184 19524 17196
rect 17267 17156 19104 17184
rect 19479 17156 19524 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 16758 17116 16764 17128
rect 14976 17088 15021 17116
rect 15672 17088 16764 17116
rect 14976 17076 14982 17088
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 15470 17048 15476 17060
rect 14108 17020 15476 17048
rect 12713 17011 12771 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16206 17008 16212 17060
rect 16264 17048 16270 17060
rect 17696 17048 17724 17079
rect 19076 17057 19104 17156
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 22035 17187 22093 17193
rect 22035 17184 22047 17187
rect 20036 17156 22047 17184
rect 20036 17144 20042 17156
rect 22035 17153 22047 17156
rect 22081 17153 22093 17187
rect 23078 17184 23106 17292
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 24728 17292 25268 17320
rect 24728 17280 24734 17292
rect 23198 17212 23204 17264
rect 23256 17252 23262 17264
rect 23256 17224 24992 17252
rect 23256 17212 23262 17224
rect 24486 17184 24492 17196
rect 23078 17156 24492 17184
rect 22035 17147 22093 17153
rect 24486 17144 24492 17156
rect 24544 17144 24550 17196
rect 24762 17144 24768 17196
rect 24820 17184 24826 17196
rect 24964 17193 24992 17224
rect 24857 17187 24915 17193
rect 24857 17184 24869 17187
rect 24820 17156 24869 17184
rect 24820 17144 24826 17156
rect 24857 17153 24869 17156
rect 24903 17153 24915 17187
rect 24857 17147 24915 17153
rect 24949 17187 25007 17193
rect 24949 17153 24961 17187
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 25038 17144 25044 17196
rect 25096 17184 25102 17196
rect 25240 17193 25268 17292
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 25961 17323 26019 17329
rect 25961 17320 25973 17323
rect 25464 17292 25973 17320
rect 25464 17280 25470 17292
rect 25961 17289 25973 17292
rect 26007 17289 26019 17323
rect 25961 17283 26019 17289
rect 25976 17252 26004 17283
rect 26050 17280 26056 17332
rect 26108 17320 26114 17332
rect 26108 17292 28120 17320
rect 26108 17280 26114 17292
rect 28092 17252 28120 17292
rect 28166 17280 28172 17332
rect 28224 17320 28230 17332
rect 28445 17323 28503 17329
rect 28445 17320 28457 17323
rect 28224 17292 28457 17320
rect 28224 17280 28230 17292
rect 28445 17289 28457 17292
rect 28491 17289 28503 17323
rect 28445 17283 28503 17289
rect 29181 17323 29239 17329
rect 29181 17289 29193 17323
rect 29227 17320 29239 17323
rect 29546 17320 29552 17332
rect 29227 17292 29552 17320
rect 29227 17289 29239 17292
rect 29181 17283 29239 17289
rect 29546 17280 29552 17292
rect 29604 17280 29610 17332
rect 30466 17320 30472 17332
rect 30116 17292 30472 17320
rect 30116 17252 30144 17292
rect 30466 17280 30472 17292
rect 30524 17320 30530 17332
rect 30834 17320 30840 17332
rect 30524 17292 30840 17320
rect 30524 17280 30530 17292
rect 30834 17280 30840 17292
rect 30892 17280 30898 17332
rect 31018 17280 31024 17332
rect 31076 17320 31082 17332
rect 31573 17323 31631 17329
rect 31573 17320 31585 17323
rect 31076 17292 31585 17320
rect 31076 17280 31082 17292
rect 31573 17289 31585 17292
rect 31619 17289 31631 17323
rect 32582 17320 32588 17332
rect 32543 17292 32588 17320
rect 31573 17283 31631 17289
rect 32582 17280 32588 17292
rect 32640 17320 32646 17332
rect 33594 17320 33600 17332
rect 32640 17292 33600 17320
rect 32640 17280 32646 17292
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 25976 17224 27200 17252
rect 25225 17187 25283 17193
rect 25096 17156 25141 17184
rect 25096 17144 25102 17156
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25271 17156 25360 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25332 17128 25360 17156
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 27172 17193 27200 17224
rect 28092 17224 30144 17252
rect 28092 17193 28120 17224
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25464 17156 25881 17184
rect 25464 17144 25470 17156
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 26973 17187 27031 17193
rect 26973 17153 26985 17187
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 28077 17187 28135 17193
rect 28077 17153 28089 17187
rect 28123 17153 28135 17187
rect 28077 17147 28135 17153
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 21726 17116 21732 17128
rect 19208 17088 21732 17116
rect 19208 17076 19214 17088
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 22278 17116 22284 17128
rect 22239 17088 22284 17116
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 22646 17076 22652 17128
rect 22704 17116 22710 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22704 17088 22753 17116
rect 22704 17076 22710 17088
rect 22741 17085 22753 17088
rect 22787 17085 22799 17119
rect 22741 17079 22799 17085
rect 25314 17076 25320 17128
rect 25372 17076 25378 17128
rect 26988 17116 27016 17147
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 30116 17193 30144 17224
rect 30392 17224 32444 17252
rect 29365 17187 29423 17193
rect 29365 17184 29377 17187
rect 29052 17156 29377 17184
rect 29052 17144 29058 17156
rect 29365 17153 29377 17156
rect 29411 17153 29423 17187
rect 29365 17147 29423 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17153 30159 17187
rect 30101 17147 30159 17153
rect 27890 17116 27896 17128
rect 26988 17088 27896 17116
rect 27890 17076 27896 17088
rect 27948 17076 27954 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17085 28227 17119
rect 28169 17079 28227 17085
rect 16264 17020 17724 17048
rect 19061 17051 19119 17057
rect 16264 17008 16270 17020
rect 19061 17017 19073 17051
rect 19107 17048 19119 17051
rect 21542 17048 21548 17060
rect 19107 17020 21548 17048
rect 19107 17017 19119 17020
rect 19061 17011 19119 17017
rect 21542 17008 21548 17020
rect 21600 17008 21606 17060
rect 24302 17008 24308 17060
rect 24360 17048 24366 17060
rect 27430 17048 27436 17060
rect 24360 17020 27436 17048
rect 24360 17008 24366 17020
rect 27430 17008 27436 17020
rect 27488 17008 27494 17060
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 28184 17048 28212 17079
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 29641 17119 29699 17125
rect 29641 17116 29653 17119
rect 28776 17088 29653 17116
rect 28776 17076 28782 17088
rect 29641 17085 29653 17088
rect 29687 17085 29699 17119
rect 30392 17116 30420 17224
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17184 30527 17187
rect 31018 17184 31024 17196
rect 30515 17156 31024 17184
rect 30515 17153 30527 17156
rect 30469 17147 30527 17153
rect 31018 17144 31024 17156
rect 31076 17184 31082 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 31076 17156 31217 17184
rect 31076 17144 31082 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 31297 17187 31355 17193
rect 31297 17153 31309 17187
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17184 31447 17187
rect 31662 17184 31668 17196
rect 31435 17156 31668 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 31312 17116 31340 17147
rect 31662 17144 31668 17156
rect 31720 17144 31726 17196
rect 32214 17184 32220 17196
rect 32175 17156 32220 17184
rect 32214 17144 32220 17156
rect 32272 17144 32278 17196
rect 32416 17193 32444 17224
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 32401 17187 32459 17193
rect 32401 17153 32413 17187
rect 32447 17184 32459 17187
rect 33318 17184 33324 17196
rect 32447 17156 33324 17184
rect 32447 17153 32459 17156
rect 32401 17147 32459 17153
rect 32232 17116 32260 17144
rect 30392 17088 30788 17116
rect 31312 17088 32260 17116
rect 29641 17079 29699 17085
rect 29178 17048 29184 17060
rect 27764 17020 29184 17048
rect 27764 17008 27770 17020
rect 29178 17008 29184 17020
rect 29236 17008 29242 17060
rect 29270 17008 29276 17060
rect 29328 17048 29334 17060
rect 29549 17051 29607 17057
rect 29549 17048 29561 17051
rect 29328 17020 29561 17048
rect 29328 17008 29334 17020
rect 29549 17017 29561 17020
rect 29595 17048 29607 17051
rect 30653 17051 30711 17057
rect 30653 17048 30665 17051
rect 29595 17020 30665 17048
rect 29595 17017 29607 17020
rect 29549 17011 29607 17017
rect 30653 17017 30665 17020
rect 30699 17017 30711 17051
rect 30653 17011 30711 17017
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12526 16980 12532 16992
rect 12487 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 14001 16983 14059 16989
rect 14001 16949 14013 16983
rect 14047 16980 14059 16983
rect 15102 16980 15108 16992
rect 14047 16952 15108 16980
rect 14047 16949 14059 16952
rect 14001 16943 14059 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 19242 16980 19248 16992
rect 17184 16952 19248 16980
rect 17184 16940 17190 16952
rect 19242 16940 19248 16952
rect 19300 16980 19306 16992
rect 20530 16980 20536 16992
rect 19300 16952 20536 16980
rect 19300 16940 19306 16952
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20809 16983 20867 16989
rect 20809 16980 20821 16983
rect 20680 16952 20821 16980
rect 20680 16940 20686 16952
rect 20809 16949 20821 16952
rect 20855 16949 20867 16983
rect 20809 16943 20867 16949
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 20956 16952 21833 16980
rect 20956 16940 20962 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 21910 16940 21916 16992
rect 21968 16980 21974 16992
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 21968 16952 22201 16980
rect 21968 16940 21974 16952
rect 22189 16949 22201 16952
rect 22235 16949 22247 16983
rect 22189 16943 22247 16949
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 24026 16980 24032 16992
rect 22980 16952 24032 16980
rect 22980 16940 22986 16952
rect 24026 16940 24032 16952
rect 24084 16980 24090 16992
rect 24121 16983 24179 16989
rect 24121 16980 24133 16983
rect 24084 16952 24133 16980
rect 24084 16940 24090 16952
rect 24121 16949 24133 16952
rect 24167 16949 24179 16983
rect 27062 16980 27068 16992
rect 27023 16952 27068 16980
rect 24121 16943 24179 16949
rect 27062 16940 27068 16952
rect 27120 16940 27126 16992
rect 28261 16983 28319 16989
rect 28261 16949 28273 16983
rect 28307 16980 28319 16983
rect 28442 16980 28448 16992
rect 28307 16952 28448 16980
rect 28307 16949 28319 16952
rect 28261 16943 28319 16949
rect 28442 16940 28448 16952
rect 28500 16980 28506 16992
rect 30377 16983 30435 16989
rect 30377 16980 30389 16983
rect 28500 16952 30389 16980
rect 28500 16940 28506 16952
rect 30377 16949 30389 16952
rect 30423 16980 30435 16983
rect 30760 16980 30788 17088
rect 30834 17008 30840 17060
rect 30892 17048 30898 17060
rect 32324 17048 32352 17147
rect 33318 17144 33324 17156
rect 33376 17144 33382 17196
rect 30892 17020 32352 17048
rect 30892 17008 30898 17020
rect 30423 16952 30788 16980
rect 30423 16949 30435 16952
rect 30377 16943 30435 16949
rect 32214 16940 32220 16992
rect 32272 16980 32278 16992
rect 33042 16980 33048 16992
rect 32272 16952 33048 16980
rect 32272 16940 32278 16952
rect 33042 16940 33048 16952
rect 33100 16940 33106 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 13722 16776 13728 16788
rect 12207 16748 13728 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 13872 16748 15025 16776
rect 13872 16736 13878 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17000 16748 18429 16776
rect 17000 16736 17006 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 19978 16776 19984 16788
rect 19939 16748 19984 16776
rect 18417 16739 18475 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20530 16736 20536 16788
rect 20588 16776 20594 16788
rect 20901 16779 20959 16785
rect 20901 16776 20913 16779
rect 20588 16748 20913 16776
rect 20588 16736 20594 16748
rect 20901 16745 20913 16748
rect 20947 16745 20959 16779
rect 20901 16739 20959 16745
rect 21453 16779 21511 16785
rect 21453 16745 21465 16779
rect 21499 16776 21511 16779
rect 23658 16776 23664 16788
rect 21499 16748 23664 16776
rect 21499 16745 21511 16748
rect 21453 16739 21511 16745
rect 23658 16736 23664 16748
rect 23716 16736 23722 16788
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 24912 16748 25912 16776
rect 24912 16736 24918 16748
rect 15746 16708 15752 16720
rect 13464 16680 15752 16708
rect 11514 16640 11520 16652
rect 11427 16612 11520 16640
rect 11514 16600 11520 16612
rect 11572 16640 11578 16652
rect 12158 16640 12164 16652
rect 11572 16612 12164 16640
rect 11572 16600 11578 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16572 10839 16575
rect 11238 16572 11244 16584
rect 10827 16544 11244 16572
rect 10827 16541 10839 16544
rect 10781 16535 10839 16541
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 12618 16572 12624 16584
rect 11379 16544 12624 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 12710 16532 12716 16584
rect 12768 16572 12774 16584
rect 12768 16544 12813 16572
rect 12768 16532 12774 16544
rect 12986 16532 12992 16584
rect 13044 16572 13050 16584
rect 13464 16572 13492 16680
rect 15746 16668 15752 16680
rect 15804 16668 15810 16720
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 19150 16708 19156 16720
rect 17267 16680 19156 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 19150 16668 19156 16680
rect 19208 16668 19214 16720
rect 20070 16668 20076 16720
rect 20128 16708 20134 16720
rect 23382 16708 23388 16720
rect 20128 16680 23388 16708
rect 20128 16668 20134 16680
rect 23382 16668 23388 16680
rect 23440 16668 23446 16720
rect 25774 16708 25780 16720
rect 25036 16680 25780 16708
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14240 16612 14565 16640
rect 14240 16600 14246 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 14553 16603 14611 16609
rect 15396 16612 16405 16640
rect 13044 16544 13492 16572
rect 13044 16532 13050 16544
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 14056 16544 14289 16572
rect 14056 16532 14062 16544
rect 14277 16541 14289 16544
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 14424 16544 14473 16572
rect 14424 16532 14430 16544
rect 14461 16541 14473 16544
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 14734 16572 14740 16584
rect 14691 16544 14740 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 12069 16507 12127 16513
rect 12069 16473 12081 16507
rect 12115 16504 12127 16507
rect 13078 16504 13084 16516
rect 12115 16476 13084 16504
rect 12115 16473 12127 16476
rect 12069 16467 12127 16473
rect 13078 16464 13084 16476
rect 13136 16464 13142 16516
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 14844 16504 14872 16535
rect 13228 16476 14872 16504
rect 13228 16464 13234 16476
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 10686 16436 10692 16448
rect 10643 16408 10692 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 15396 16436 15424 16612
rect 16393 16609 16405 16612
rect 16439 16640 16451 16643
rect 17126 16640 17132 16652
rect 16439 16612 17132 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17420 16612 17969 16640
rect 15654 16572 15660 16584
rect 15615 16544 15660 16572
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 15804 16544 16865 16572
rect 15804 16532 15810 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17420 16572 17448 16612
rect 17957 16609 17969 16612
rect 18003 16640 18015 16643
rect 18003 16612 18368 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 17083 16544 17448 16572
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17644 16544 17693 16572
rect 17644 16532 17650 16544
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17862 16572 17868 16584
rect 17823 16544 17868 16572
rect 17681 16535 17739 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18138 16572 18144 16584
rect 18095 16544 18144 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18340 16572 18368 16612
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 18656 16612 19625 16640
rect 18656 16600 18662 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 20714 16640 20720 16652
rect 20675 16612 20720 16640
rect 19613 16603 19671 16609
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 21450 16600 21456 16652
rect 21508 16640 21514 16652
rect 21913 16643 21971 16649
rect 21913 16640 21925 16643
rect 21508 16612 21925 16640
rect 21508 16600 21514 16612
rect 21913 16609 21925 16612
rect 21959 16609 21971 16643
rect 24302 16640 24308 16652
rect 21913 16603 21971 16609
rect 23078 16612 24308 16640
rect 18782 16572 18788 16584
rect 18340 16544 18788 16572
rect 18233 16535 18291 16541
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 16942 16504 16948 16516
rect 16255 16476 16948 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 13504 16408 15424 16436
rect 15473 16439 15531 16445
rect 13504 16396 13510 16408
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 16224 16436 16252 16467
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17402 16464 17408 16516
rect 17460 16504 17466 16516
rect 18248 16504 18276 16535
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18892 16544 19257 16572
rect 17460 16476 18276 16504
rect 17460 16464 17466 16476
rect 15519 16408 16252 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 17126 16396 17132 16448
rect 17184 16436 17190 16448
rect 17586 16436 17592 16448
rect 17184 16408 17592 16436
rect 17184 16396 17190 16408
rect 17586 16396 17592 16408
rect 17644 16436 17650 16448
rect 18892 16436 18920 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 19444 16504 19472 16535
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 19797 16575 19855 16581
rect 19576 16544 19621 16572
rect 19576 16532 19582 16544
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 19208 16476 19472 16504
rect 19208 16464 19214 16476
rect 17644 16408 18920 16436
rect 19812 16436 19840 16535
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 20496 16544 20637 16572
rect 20496 16532 20502 16544
rect 20625 16541 20637 16544
rect 20671 16572 20683 16575
rect 20671 16544 21496 16572
rect 20671 16541 20683 16544
rect 20625 16535 20683 16541
rect 20990 16464 20996 16516
rect 21048 16504 21054 16516
rect 21468 16504 21496 16544
rect 21542 16532 21548 16584
rect 21600 16572 21606 16584
rect 21637 16575 21695 16581
rect 21637 16572 21649 16575
rect 21600 16544 21649 16572
rect 21600 16532 21606 16544
rect 21637 16541 21649 16544
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 21836 16504 21864 16535
rect 22922 16532 22928 16584
rect 22980 16572 22986 16584
rect 23078 16581 23106 16612
rect 24302 16600 24308 16612
rect 24360 16600 24366 16652
rect 23063 16575 23121 16581
rect 23063 16572 23075 16575
rect 22980 16544 23075 16572
rect 22980 16532 22986 16544
rect 23063 16541 23075 16544
rect 23109 16541 23121 16575
rect 23198 16572 23204 16584
rect 23159 16544 23204 16572
rect 23063 16535 23121 16541
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 23290 16532 23296 16584
rect 23348 16572 23354 16584
rect 23477 16575 23535 16581
rect 23348 16544 23393 16572
rect 23348 16532 23354 16544
rect 23477 16541 23489 16575
rect 23523 16572 23535 16575
rect 23566 16572 23572 16584
rect 23523 16544 23572 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 25036 16581 25064 16680
rect 25774 16668 25780 16680
rect 25832 16668 25838 16720
rect 25682 16640 25688 16652
rect 25148 16612 25688 16640
rect 25148 16581 25176 16612
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 25884 16649 25912 16748
rect 26786 16736 26792 16788
rect 26844 16776 26850 16788
rect 28537 16779 28595 16785
rect 28537 16776 28549 16779
rect 26844 16748 28549 16776
rect 26844 16736 26850 16748
rect 28537 16745 28549 16748
rect 28583 16776 28595 16779
rect 29546 16776 29552 16788
rect 28583 16748 29552 16776
rect 28583 16745 28595 16748
rect 28537 16739 28595 16745
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 30285 16779 30343 16785
rect 30285 16745 30297 16779
rect 30331 16776 30343 16779
rect 30466 16776 30472 16788
rect 30331 16748 30472 16776
rect 30331 16745 30343 16748
rect 30285 16739 30343 16745
rect 30466 16736 30472 16748
rect 30524 16736 30530 16788
rect 33410 16736 33416 16788
rect 33468 16776 33474 16788
rect 33965 16779 34023 16785
rect 33965 16776 33977 16779
rect 33468 16748 33977 16776
rect 33468 16736 33474 16748
rect 33965 16745 33977 16748
rect 34011 16745 34023 16779
rect 33965 16739 34023 16745
rect 27249 16711 27307 16717
rect 27249 16677 27261 16711
rect 27295 16708 27307 16711
rect 27430 16708 27436 16720
rect 27295 16680 27436 16708
rect 27295 16677 27307 16680
rect 27249 16671 27307 16677
rect 27430 16668 27436 16680
rect 27488 16668 27494 16720
rect 29178 16668 29184 16720
rect 29236 16708 29242 16720
rect 30834 16708 30840 16720
rect 29236 16680 30840 16708
rect 29236 16668 29242 16680
rect 30834 16668 30840 16680
rect 30892 16668 30898 16720
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16609 25927 16643
rect 29730 16640 29736 16652
rect 25869 16603 25927 16609
rect 27908 16612 29736 16640
rect 25021 16575 25079 16581
rect 25021 16541 25033 16575
rect 25067 16541 25079 16575
rect 25021 16535 25079 16541
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 25409 16575 25467 16581
rect 25280 16544 25325 16572
rect 25280 16532 25286 16544
rect 25409 16541 25421 16575
rect 25455 16572 25467 16575
rect 25590 16572 25596 16584
rect 25455 16544 25596 16572
rect 25455 16541 25467 16544
rect 25409 16535 25467 16541
rect 25590 16532 25596 16544
rect 25648 16572 25654 16584
rect 27709 16575 27767 16581
rect 25648 16544 27660 16572
rect 25648 16532 25654 16544
rect 21048 16476 21093 16504
rect 21468 16476 21864 16504
rect 22833 16507 22891 16513
rect 21048 16464 21054 16476
rect 22833 16473 22845 16507
rect 22879 16504 22891 16507
rect 26114 16507 26172 16513
rect 26114 16504 26126 16507
rect 22879 16476 26126 16504
rect 22879 16473 22891 16476
rect 22833 16467 22891 16473
rect 26114 16473 26126 16476
rect 26160 16473 26172 16507
rect 27632 16504 27660 16544
rect 27709 16541 27721 16575
rect 27755 16572 27767 16575
rect 27798 16572 27804 16584
rect 27755 16544 27804 16572
rect 27755 16541 27767 16544
rect 27709 16535 27767 16541
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 27908 16581 27936 16612
rect 29730 16600 29736 16612
rect 29788 16600 29794 16652
rect 31389 16643 31447 16649
rect 31389 16609 31401 16643
rect 31435 16640 31447 16643
rect 32214 16640 32220 16652
rect 31435 16612 32220 16640
rect 31435 16609 31447 16612
rect 31389 16603 31447 16609
rect 32214 16600 32220 16612
rect 32272 16600 32278 16652
rect 32861 16643 32919 16649
rect 32324 16612 32536 16640
rect 27893 16575 27951 16581
rect 27893 16541 27905 16575
rect 27939 16541 27951 16575
rect 27893 16535 27951 16541
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16572 28503 16575
rect 30374 16572 30380 16584
rect 28491 16544 30380 16572
rect 28491 16541 28503 16544
rect 28445 16535 28503 16541
rect 30374 16532 30380 16544
rect 30432 16532 30438 16584
rect 31113 16575 31171 16581
rect 31113 16541 31125 16575
rect 31159 16541 31171 16575
rect 31113 16535 31171 16541
rect 28350 16504 28356 16516
rect 27632 16476 28356 16504
rect 26114 16467 26172 16473
rect 28350 16464 28356 16476
rect 28408 16464 28414 16516
rect 30193 16507 30251 16513
rect 30193 16473 30205 16507
rect 30239 16504 30251 16507
rect 30466 16504 30472 16516
rect 30239 16476 30472 16504
rect 30239 16473 30251 16476
rect 30193 16467 30251 16473
rect 30466 16464 30472 16476
rect 30524 16504 30530 16516
rect 31128 16504 31156 16535
rect 31662 16532 31668 16584
rect 31720 16572 31726 16584
rect 32324 16572 32352 16612
rect 31720 16544 32352 16572
rect 32401 16575 32459 16581
rect 31720 16532 31726 16544
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32508 16572 32536 16612
rect 32861 16609 32873 16643
rect 32907 16640 32919 16643
rect 33134 16640 33140 16652
rect 32907 16612 33140 16640
rect 32907 16609 32919 16612
rect 32861 16603 32919 16609
rect 33134 16600 33140 16612
rect 33192 16600 33198 16652
rect 33520 16612 33824 16640
rect 32769 16575 32827 16581
rect 32769 16572 32781 16575
rect 32508 16544 32781 16572
rect 32401 16535 32459 16541
rect 32769 16541 32781 16544
rect 32815 16541 32827 16575
rect 32950 16572 32956 16584
rect 32911 16544 32956 16572
rect 32769 16535 32827 16541
rect 30524 16476 31156 16504
rect 30524 16464 30530 16476
rect 21358 16436 21364 16448
rect 19812 16408 21364 16436
rect 17644 16396 17650 16408
rect 21358 16396 21364 16408
rect 21416 16396 21422 16448
rect 24765 16439 24823 16445
rect 24765 16405 24777 16439
rect 24811 16436 24823 16439
rect 25590 16436 25596 16448
rect 24811 16408 25596 16436
rect 24811 16405 24823 16408
rect 24765 16399 24823 16405
rect 25590 16396 25596 16408
rect 25648 16396 25654 16448
rect 27893 16439 27951 16445
rect 27893 16405 27905 16439
rect 27939 16436 27951 16439
rect 28166 16436 28172 16448
rect 27939 16408 28172 16436
rect 27939 16405 27951 16408
rect 27893 16399 27951 16405
rect 28166 16396 28172 16408
rect 28224 16396 28230 16448
rect 32122 16396 32128 16448
rect 32180 16436 32186 16448
rect 32416 16436 32444 16535
rect 32784 16504 32812 16535
rect 32950 16532 32956 16544
rect 33008 16572 33014 16584
rect 33520 16572 33548 16612
rect 33796 16581 33824 16612
rect 33008 16544 33548 16572
rect 33597 16575 33655 16581
rect 33008 16532 33014 16544
rect 33597 16541 33609 16575
rect 33643 16541 33655 16575
rect 33597 16535 33655 16541
rect 33689 16575 33747 16581
rect 33689 16541 33701 16575
rect 33735 16541 33747 16575
rect 33689 16535 33747 16541
rect 33781 16575 33839 16581
rect 33781 16541 33793 16575
rect 33827 16574 33839 16575
rect 33827 16546 33861 16574
rect 33827 16541 33839 16546
rect 33781 16535 33839 16541
rect 33612 16504 33640 16535
rect 32784 16476 33640 16504
rect 33704 16436 33732 16535
rect 32180 16408 33732 16436
rect 32180 16396 32186 16408
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 15654 16232 15660 16244
rect 13136 16204 13676 16232
rect 13136 16192 13142 16204
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16164 13415 16167
rect 13446 16164 13452 16176
rect 13403 16136 13452 16164
rect 13403 16133 13415 16136
rect 13357 16127 13415 16133
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 13538 16124 13544 16176
rect 13596 16173 13602 16176
rect 13596 16167 13615 16173
rect 13603 16133 13615 16167
rect 13648 16164 13676 16204
rect 14568 16204 15660 16232
rect 14568 16176 14596 16204
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 17862 16232 17868 16244
rect 16816 16204 17868 16232
rect 16816 16192 16822 16204
rect 17862 16192 17868 16204
rect 17920 16232 17926 16244
rect 19150 16232 19156 16244
rect 17920 16204 19156 16232
rect 17920 16192 17926 16204
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 22189 16235 22247 16241
rect 21600 16204 22048 16232
rect 21600 16192 21606 16204
rect 14550 16164 14556 16176
rect 13648 16136 14556 16164
rect 13596 16127 13615 16133
rect 13596 16124 13602 16127
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 14660 16136 16988 16164
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 11698 16096 11704 16108
rect 10459 16068 11704 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12710 16096 12716 16108
rect 12207 16068 12434 16096
rect 12623 16068 12716 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12406 15960 12434 16068
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 13556 16096 13584 16124
rect 14458 16096 14464 16108
rect 12943 16068 13584 16096
rect 14419 16068 14464 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14660 16105 14688 16136
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14568 16068 14657 16096
rect 12728 16028 12756 16056
rect 13630 16028 13636 16040
rect 12728 16000 13636 16028
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 14366 15988 14372 16040
rect 14424 16028 14430 16040
rect 14568 16028 14596 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15243 16068 15853 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 14734 16028 14740 16040
rect 14424 16000 14596 16028
rect 14695 16000 14740 16028
rect 14424 15988 14430 16000
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 14826 15988 14832 16040
rect 14884 16028 14890 16040
rect 14884 16000 14929 16028
rect 14884 15988 14890 16000
rect 13725 15963 13783 15969
rect 13725 15960 13737 15963
rect 12406 15932 13737 15960
rect 13725 15929 13737 15932
rect 13771 15929 13783 15963
rect 13725 15923 13783 15929
rect 14274 15920 14280 15972
rect 14332 15960 14338 15972
rect 15028 15960 15056 16059
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16669 16099 16727 16105
rect 15988 16068 16252 16096
rect 15988 16056 15994 16068
rect 16114 16028 16120 16040
rect 16075 16000 16120 16028
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16224 16028 16252 16068
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 16758 16096 16764 16108
rect 16715 16068 16764 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 16960 16105 16988 16136
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 19702 16164 19708 16176
rect 18012 16136 19708 16164
rect 18012 16124 18018 16136
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 22020 16173 22048 16204
rect 22189 16201 22201 16235
rect 22235 16232 22247 16235
rect 23290 16232 23296 16244
rect 22235 16204 23296 16232
rect 22235 16201 22247 16204
rect 22189 16195 22247 16201
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 26329 16235 26387 16241
rect 26329 16232 26341 16235
rect 25280 16204 26341 16232
rect 25280 16192 25286 16204
rect 26329 16201 26341 16204
rect 26375 16201 26387 16235
rect 30282 16232 30288 16244
rect 30243 16204 30288 16232
rect 26329 16195 26387 16201
rect 30282 16192 30288 16204
rect 30340 16192 30346 16244
rect 32398 16192 32404 16244
rect 32456 16232 32462 16244
rect 32677 16235 32735 16241
rect 32677 16232 32689 16235
rect 32456 16204 32689 16232
rect 32456 16192 32462 16204
rect 32677 16201 32689 16204
rect 32723 16201 32735 16235
rect 33318 16232 33324 16244
rect 33279 16204 33324 16232
rect 32677 16195 32735 16201
rect 33318 16192 33324 16204
rect 33376 16192 33382 16244
rect 22005 16167 22063 16173
rect 19904 16136 21956 16164
rect 19904 16108 19932 16136
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17678 16096 17684 16108
rect 16991 16068 17684 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 18598 16096 18604 16108
rect 17788 16068 18460 16096
rect 18559 16068 18604 16096
rect 17788 16028 17816 16068
rect 16224 16000 17816 16028
rect 18230 15988 18236 16040
rect 18288 16028 18294 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18288 16000 18337 16028
rect 18288 15988 18294 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18432 16028 18460 16068
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 19886 16096 19892 16108
rect 19843 16068 19892 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 20070 16105 20076 16108
rect 20064 16059 20076 16105
rect 20128 16096 20134 16108
rect 20128 16068 20164 16096
rect 20070 16056 20076 16059
rect 20128 16056 20134 16068
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21692 16068 21833 16096
rect 21692 16056 21698 16068
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 21928 16096 21956 16136
rect 22005 16133 22017 16167
rect 22051 16133 22063 16167
rect 24854 16164 24860 16176
rect 22005 16127 22063 16133
rect 24136 16136 24860 16164
rect 22646 16096 22652 16108
rect 21928 16068 22652 16096
rect 21821 16059 21879 16065
rect 19610 16028 19616 16040
rect 18432 16000 19616 16028
rect 18325 15991 18383 15997
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 14332 15932 15056 15960
rect 14332 15920 14338 15932
rect 15102 15920 15108 15972
rect 15160 15960 15166 15972
rect 16132 15960 16160 15988
rect 19794 15960 19800 15972
rect 15160 15932 15792 15960
rect 16132 15932 19800 15960
rect 15160 15920 15166 15932
rect 15764 15904 15792 15932
rect 19794 15920 19800 15932
rect 19852 15920 19858 15972
rect 20990 15960 20996 15972
rect 20732 15932 20996 15960
rect 10226 15892 10232 15904
rect 10187 15864 10232 15892
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 11977 15895 12035 15901
rect 11977 15861 11989 15895
rect 12023 15892 12035 15895
rect 12250 15892 12256 15904
rect 12023 15864 12256 15892
rect 12023 15861 12035 15864
rect 11977 15855 12035 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 13538 15892 13544 15904
rect 13499 15864 13544 15892
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15344 15864 15669 15892
rect 15344 15852 15350 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15804 15864 16037 15892
rect 15804 15852 15810 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 18230 15852 18236 15904
rect 18288 15892 18294 15904
rect 20732 15892 20760 15932
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 21836 15960 21864 16059
rect 22646 16056 22652 16068
rect 22704 16096 22710 16108
rect 24136 16105 24164 16136
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 26145 16167 26203 16173
rect 26145 16164 26157 16167
rect 25004 16136 26157 16164
rect 25004 16124 25010 16136
rect 26145 16133 26157 16136
rect 26191 16133 26203 16167
rect 26145 16127 26203 16133
rect 24394 16105 24400 16108
rect 24121 16099 24179 16105
rect 24121 16096 24133 16099
rect 22704 16068 24133 16096
rect 22704 16056 22710 16068
rect 24121 16065 24133 16068
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 24388 16059 24400 16105
rect 24452 16096 24458 16108
rect 25961 16099 26019 16105
rect 24452 16068 24488 16096
rect 24394 16056 24400 16059
rect 24452 16056 24458 16068
rect 25961 16065 25973 16099
rect 26007 16096 26019 16099
rect 26970 16096 26976 16108
rect 26007 16068 26976 16096
rect 26007 16065 26019 16068
rect 25961 16059 26019 16065
rect 22833 16031 22891 16037
rect 22833 15997 22845 16031
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 23109 16031 23167 16037
rect 23109 15997 23121 16031
rect 23155 16028 23167 16031
rect 23198 16028 23204 16040
rect 23155 16000 23204 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 22002 15960 22008 15972
rect 21836 15932 22008 15960
rect 22002 15920 22008 15932
rect 22060 15960 22066 15972
rect 22848 15960 22876 15991
rect 23198 15988 23204 16000
rect 23256 15988 23262 16040
rect 23566 15960 23572 15972
rect 22060 15932 22324 15960
rect 22848 15932 23572 15960
rect 22060 15920 22066 15932
rect 18288 15864 20760 15892
rect 18288 15852 18294 15864
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21177 15895 21235 15901
rect 21177 15892 21189 15895
rect 20864 15864 21189 15892
rect 20864 15852 20870 15864
rect 21177 15861 21189 15864
rect 21223 15861 21235 15895
rect 21177 15855 21235 15861
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22186 15892 22192 15904
rect 21968 15864 22192 15892
rect 21968 15852 21974 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22296 15892 22324 15932
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 25976 15960 26004 16059
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 27065 16099 27123 16105
rect 27065 16065 27077 16099
rect 27111 16096 27123 16099
rect 27706 16096 27712 16108
rect 27111 16068 27712 16096
rect 27111 16065 27123 16068
rect 27065 16059 27123 16065
rect 27706 16056 27712 16068
rect 27764 16056 27770 16108
rect 27982 16096 27988 16108
rect 27943 16068 27988 16096
rect 27982 16056 27988 16068
rect 28040 16056 28046 16108
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16065 28135 16099
rect 28077 16059 28135 16065
rect 27890 15988 27896 16040
rect 27948 16028 27954 16040
rect 28092 16028 28120 16059
rect 28166 16056 28172 16108
rect 28224 16096 28230 16108
rect 28350 16096 28356 16108
rect 28224 16068 28269 16096
rect 28311 16068 28356 16096
rect 28224 16056 28230 16068
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28442 16056 28448 16108
rect 28500 16096 28506 16108
rect 28813 16099 28871 16105
rect 28813 16096 28825 16099
rect 28500 16068 28825 16096
rect 28500 16056 28506 16068
rect 28813 16065 28825 16068
rect 28859 16065 28871 16099
rect 28813 16059 28871 16065
rect 29733 16099 29791 16105
rect 29733 16065 29745 16099
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 30101 16099 30159 16105
rect 30101 16065 30113 16099
rect 30147 16096 30159 16099
rect 30745 16099 30803 16105
rect 30745 16096 30757 16099
rect 30147 16068 30757 16096
rect 30147 16065 30159 16068
rect 30101 16059 30159 16065
rect 30745 16065 30757 16068
rect 30791 16096 30803 16099
rect 31202 16096 31208 16108
rect 30791 16068 31208 16096
rect 30791 16065 30803 16068
rect 30745 16059 30803 16065
rect 27948 16000 28120 16028
rect 29748 16028 29776 16059
rect 31202 16056 31208 16068
rect 31260 16056 31266 16108
rect 32122 16096 32128 16108
rect 31312 16068 32128 16096
rect 30650 16028 30656 16040
rect 29748 16000 30656 16028
rect 27948 15988 27954 16000
rect 30650 15988 30656 16000
rect 30708 15988 30714 16040
rect 31018 16028 31024 16040
rect 30979 16000 31024 16028
rect 31018 15988 31024 16000
rect 31076 16028 31082 16040
rect 31312 16028 31340 16068
rect 32122 16056 32128 16068
rect 32180 16056 32186 16108
rect 33229 16099 33287 16105
rect 33229 16065 33241 16099
rect 33275 16065 33287 16099
rect 33229 16059 33287 16065
rect 31076 16000 31340 16028
rect 31076 15988 31082 16000
rect 31662 15988 31668 16040
rect 31720 16028 31726 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 31720 16000 32413 16028
rect 31720 15988 31726 16000
rect 32401 15997 32413 16000
rect 32447 16028 32459 16031
rect 33244 16028 33272 16059
rect 32447 16000 33272 16028
rect 32447 15997 32459 16000
rect 32401 15991 32459 15997
rect 25056 15932 26004 15960
rect 27157 15963 27215 15969
rect 25056 15892 25084 15932
rect 27157 15929 27169 15963
rect 27203 15960 27215 15963
rect 28534 15960 28540 15972
rect 27203 15932 28540 15960
rect 27203 15929 27215 15932
rect 27157 15923 27215 15929
rect 28534 15920 28540 15932
rect 28592 15960 28598 15972
rect 28718 15960 28724 15972
rect 28592 15932 28724 15960
rect 28592 15920 28598 15932
rect 28718 15920 28724 15932
rect 28776 15920 28782 15972
rect 30466 15960 30472 15972
rect 30116 15932 30472 15960
rect 22296 15864 25084 15892
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 25501 15895 25559 15901
rect 25501 15892 25513 15895
rect 25464 15864 25513 15892
rect 25464 15852 25470 15864
rect 25501 15861 25513 15864
rect 25547 15861 25559 15895
rect 25501 15855 25559 15861
rect 27709 15895 27767 15901
rect 27709 15861 27721 15895
rect 27755 15892 27767 15895
rect 28810 15892 28816 15904
rect 27755 15864 28816 15892
rect 27755 15861 27767 15864
rect 27709 15855 27767 15861
rect 28810 15852 28816 15864
rect 28868 15852 28874 15904
rect 28902 15852 28908 15904
rect 28960 15892 28966 15904
rect 30116 15901 30144 15932
rect 30466 15920 30472 15932
rect 30524 15920 30530 15972
rect 30101 15895 30159 15901
rect 28960 15864 29005 15892
rect 28960 15852 28966 15864
rect 30101 15861 30113 15895
rect 30147 15861 30159 15895
rect 30101 15855 30159 15861
rect 32493 15895 32551 15901
rect 32493 15861 32505 15895
rect 32539 15892 32551 15895
rect 32950 15892 32956 15904
rect 32539 15864 32956 15892
rect 32539 15861 32551 15864
rect 32493 15855 32551 15861
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 16540 15660 18521 15688
rect 16540 15648 16546 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 24394 15688 24400 15700
rect 24355 15660 24400 15688
rect 18509 15651 18567 15657
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 27062 15688 27068 15700
rect 24971 15660 27068 15688
rect 10873 15623 10931 15629
rect 10873 15589 10885 15623
rect 10919 15620 10931 15623
rect 11790 15620 11796 15632
rect 10919 15592 11796 15620
rect 10919 15589 10931 15592
rect 10873 15583 10931 15589
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 14826 15580 14832 15632
rect 14884 15620 14890 15632
rect 16390 15620 16396 15632
rect 14884 15592 16396 15620
rect 14884 15580 14890 15592
rect 10502 15512 10508 15564
rect 10560 15552 10566 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 10560 15524 11713 15552
rect 10560 15512 10566 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 14366 15512 14372 15564
rect 14424 15552 14430 15564
rect 15028 15561 15056 15592
rect 16390 15580 16396 15592
rect 16448 15580 16454 15632
rect 16574 15580 16580 15632
rect 16632 15620 16638 15632
rect 16632 15592 17356 15620
rect 16632 15580 16638 15592
rect 15013 15555 15071 15561
rect 14424 15524 14872 15552
rect 14424 15512 14430 15524
rect 9490 15484 9496 15496
rect 9403 15456 9496 15484
rect 9490 15444 9496 15456
rect 9548 15484 9554 15496
rect 12158 15484 12164 15496
rect 9548 15456 12164 15484
rect 9548 15444 9554 15456
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12417 15487 12475 15493
rect 12417 15484 12429 15487
rect 12308 15456 12429 15484
rect 12308 15444 12314 15456
rect 12417 15453 12429 15456
rect 12463 15453 12475 15487
rect 12417 15447 12475 15453
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 14844 15493 14872 15524
rect 15013 15521 15025 15555
rect 15059 15521 15071 15555
rect 15930 15552 15936 15564
rect 15013 15515 15071 15521
rect 15120 15524 15936 15552
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14516 15456 14657 15484
rect 14516 15444 14522 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15484 14979 15487
rect 15120 15484 15148 15524
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15552 16359 15555
rect 16758 15552 16764 15564
rect 16347 15524 16764 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 17328 15561 17356 15592
rect 20254 15580 20260 15632
rect 20312 15620 20318 15632
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 20312 15592 21189 15620
rect 20312 15580 20318 15592
rect 21177 15589 21189 15592
rect 21223 15589 21235 15623
rect 21818 15620 21824 15632
rect 21177 15583 21235 15589
rect 21744 15592 21824 15620
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 17000 15524 17049 15552
rect 17000 15512 17006 15524
rect 17037 15521 17049 15524
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15552 17371 15555
rect 17954 15552 17960 15564
rect 17359 15524 17960 15552
rect 17359 15521 17371 15524
rect 17313 15515 17371 15521
rect 14967 15456 15148 15484
rect 15197 15487 15255 15493
rect 14967 15453 14979 15456
rect 14921 15447 14979 15453
rect 15197 15453 15209 15487
rect 15243 15484 15255 15487
rect 15838 15484 15844 15496
rect 15243 15456 15844 15484
rect 15243 15453 15255 15456
rect 15197 15447 15255 15453
rect 9760 15419 9818 15425
rect 9760 15385 9772 15419
rect 9806 15385 9818 15419
rect 11330 15416 11336 15428
rect 11291 15388 11336 15416
rect 9760 15379 9818 15385
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 9784 15348 9812 15379
rect 11330 15376 11336 15388
rect 11388 15376 11394 15428
rect 11517 15419 11575 15425
rect 11517 15385 11529 15419
rect 11563 15385 11575 15419
rect 14660 15416 14688 15447
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16209 15447 16267 15453
rect 16040 15416 16068 15447
rect 14660 15388 16068 15416
rect 16224 15416 16252 15447
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16666 15484 16672 15496
rect 16623 15456 16672 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 17052 15484 17080 15515
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 19242 15552 19248 15564
rect 19203 15524 19248 15552
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 20990 15552 20996 15564
rect 19852 15524 20996 15552
rect 19852 15512 19858 15524
rect 20990 15512 20996 15524
rect 21048 15552 21054 15564
rect 21744 15561 21772 15592
rect 21818 15580 21824 15592
rect 21876 15580 21882 15632
rect 22830 15580 22836 15632
rect 22888 15620 22894 15632
rect 24762 15620 24768 15632
rect 22888 15592 24768 15620
rect 22888 15580 22894 15592
rect 24762 15580 24768 15592
rect 24820 15580 24826 15632
rect 21637 15555 21695 15561
rect 21637 15552 21649 15555
rect 21048 15524 21649 15552
rect 21048 15512 21054 15524
rect 21637 15521 21649 15524
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15521 21787 15555
rect 24578 15552 24584 15564
rect 21729 15515 21787 15521
rect 22940 15524 24584 15552
rect 18138 15484 18144 15496
rect 17052 15456 18144 15484
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15484 18291 15487
rect 18506 15484 18512 15496
rect 18279 15456 18512 15484
rect 18279 15453 18291 15456
rect 18233 15447 18291 15453
rect 18506 15444 18512 15456
rect 18564 15484 18570 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18564 15456 18705 15484
rect 18564 15444 18570 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15484 19579 15487
rect 20254 15484 20260 15496
rect 19567 15456 20260 15484
rect 19567 15453 19579 15456
rect 19521 15447 19579 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20533 15487 20591 15493
rect 20533 15453 20545 15487
rect 20579 15484 20591 15487
rect 21450 15484 21456 15496
rect 20579 15456 21456 15484
rect 20579 15453 20591 15456
rect 20533 15447 20591 15453
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 21818 15444 21824 15496
rect 21876 15484 21882 15496
rect 22940 15493 22968 15524
rect 24578 15512 24584 15524
rect 24636 15552 24642 15564
rect 24636 15524 24808 15552
rect 24636 15512 24642 15524
rect 22649 15487 22707 15493
rect 22649 15484 22661 15487
rect 21876 15456 22661 15484
rect 21876 15444 21882 15456
rect 22649 15453 22661 15456
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 24670 15484 24676 15496
rect 24631 15456 24676 15484
rect 22925 15447 22983 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 24780 15493 24808 15524
rect 24762 15487 24820 15493
rect 24762 15453 24774 15487
rect 24808 15453 24820 15487
rect 24762 15447 24820 15453
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15484 24915 15487
rect 24971 15484 24999 15660
rect 27062 15648 27068 15660
rect 27120 15648 27126 15700
rect 30466 15648 30472 15700
rect 30524 15688 30530 15700
rect 30929 15691 30987 15697
rect 30929 15688 30941 15691
rect 30524 15660 30941 15688
rect 30524 15648 30530 15660
rect 30929 15657 30941 15660
rect 30975 15657 30987 15691
rect 30929 15651 30987 15657
rect 25038 15580 25044 15632
rect 25096 15580 25102 15632
rect 26878 15620 26884 15632
rect 26839 15592 26884 15620
rect 26878 15580 26884 15592
rect 26936 15580 26942 15632
rect 25056 15552 25084 15580
rect 25501 15555 25559 15561
rect 25501 15552 25513 15555
rect 25056 15524 25513 15552
rect 25501 15521 25513 15524
rect 25547 15521 25559 15555
rect 25501 15515 25559 15521
rect 28350 15512 28356 15564
rect 28408 15552 28414 15564
rect 28408 15524 28488 15552
rect 28408 15512 28414 15524
rect 24903 15456 24999 15484
rect 25041 15487 25099 15493
rect 24903 15453 24915 15456
rect 24857 15447 24915 15453
rect 25041 15453 25053 15487
rect 25087 15484 25099 15487
rect 25314 15484 25320 15496
rect 25087 15456 25320 15484
rect 25087 15453 25099 15456
rect 25041 15447 25099 15453
rect 25314 15444 25320 15456
rect 25372 15444 25378 15496
rect 25590 15444 25596 15496
rect 25648 15484 25654 15496
rect 25757 15487 25815 15493
rect 25757 15484 25769 15487
rect 25648 15456 25769 15484
rect 25648 15444 25654 15456
rect 25757 15453 25769 15456
rect 25803 15453 25815 15487
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 25757 15447 25815 15453
rect 25884 15456 28089 15484
rect 17126 15416 17132 15428
rect 16224 15388 17132 15416
rect 11517 15379 11575 15385
rect 9732 15320 9812 15348
rect 9732 15308 9738 15320
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 11532 15348 11560 15379
rect 11020 15320 11560 15348
rect 11020 15308 11026 15320
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15381 15351 15439 15357
rect 15381 15348 15393 15351
rect 15252 15320 15393 15348
rect 15252 15308 15258 15320
rect 15381 15317 15393 15320
rect 15427 15317 15439 15351
rect 16040 15348 16068 15388
rect 17126 15376 17132 15388
rect 17184 15376 17190 15428
rect 20625 15419 20683 15425
rect 20625 15385 20637 15419
rect 20671 15416 20683 15419
rect 20714 15416 20720 15428
rect 20671 15388 20720 15416
rect 20671 15385 20683 15388
rect 20625 15379 20683 15385
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 25884 15416 25912 15456
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 27890 15416 27896 15428
rect 21468 15388 25912 15416
rect 27724 15388 27896 15416
rect 16574 15348 16580 15360
rect 16040 15320 16580 15348
rect 15381 15311 15439 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 16761 15351 16819 15357
rect 16761 15317 16773 15351
rect 16807 15348 16819 15351
rect 16850 15348 16856 15360
rect 16807 15320 16856 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 21468 15348 21496 15388
rect 17552 15320 21496 15348
rect 21545 15351 21603 15357
rect 17552 15308 17558 15320
rect 21545 15317 21557 15351
rect 21591 15348 21603 15351
rect 22462 15348 22468 15360
rect 21591 15320 22468 15348
rect 21591 15317 21603 15320
rect 21545 15311 21603 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 24578 15308 24584 15360
rect 24636 15348 24642 15360
rect 27724 15348 27752 15388
rect 27890 15376 27896 15388
rect 27948 15416 27954 15428
rect 28184 15416 28212 15447
rect 28258 15444 28264 15496
rect 28316 15484 28322 15496
rect 28460 15493 28488 15524
rect 29270 15512 29276 15564
rect 29328 15552 29334 15564
rect 29546 15552 29552 15564
rect 29328 15524 29552 15552
rect 29328 15512 29334 15524
rect 29546 15512 29552 15524
rect 29604 15512 29610 15564
rect 31662 15552 31668 15564
rect 31623 15524 31668 15552
rect 31662 15512 31668 15524
rect 31720 15512 31726 15564
rect 28445 15487 28503 15493
rect 28316 15456 28361 15484
rect 28316 15444 28322 15456
rect 28445 15453 28457 15487
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 28810 15444 28816 15496
rect 28868 15484 28874 15496
rect 29805 15487 29863 15493
rect 29805 15484 29817 15487
rect 28868 15456 29817 15484
rect 28868 15444 28874 15456
rect 29805 15453 29817 15456
rect 29851 15453 29863 15487
rect 29805 15447 29863 15453
rect 30650 15444 30656 15496
rect 30708 15484 30714 15496
rect 31389 15487 31447 15493
rect 31389 15484 31401 15487
rect 30708 15456 31401 15484
rect 30708 15444 30714 15456
rect 31389 15453 31401 15456
rect 31435 15453 31447 15487
rect 31389 15447 31447 15453
rect 27948 15388 28212 15416
rect 27948 15376 27954 15388
rect 24636 15320 27752 15348
rect 27801 15351 27859 15357
rect 24636 15308 24642 15320
rect 27801 15317 27813 15351
rect 27847 15348 27859 15351
rect 29362 15348 29368 15360
rect 27847 15320 29368 15348
rect 27847 15317 27859 15320
rect 27801 15311 27859 15317
rect 29362 15308 29368 15320
rect 29420 15308 29426 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 8849 15147 8907 15153
rect 8849 15113 8861 15147
rect 8895 15144 8907 15147
rect 9674 15144 9680 15156
rect 8895 15116 9680 15144
rect 8895 15113 8907 15116
rect 8849 15107 8907 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 21542 15144 21548 15156
rect 13504 15116 21548 15144
rect 13504 15104 13510 15116
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 22002 15144 22008 15156
rect 21867 15116 22008 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 22002 15104 22008 15116
rect 22060 15104 22066 15156
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 25590 15144 25596 15156
rect 23624 15116 25596 15144
rect 23624 15104 23630 15116
rect 9760 15079 9818 15085
rect 9048 15048 9720 15076
rect 9048 15017 9076 15048
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 14977 9091 15011
rect 9490 15008 9496 15020
rect 9451 14980 9496 15008
rect 9033 14971 9091 14977
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 9692 15008 9720 15048
rect 9760 15045 9772 15079
rect 9806 15076 9818 15079
rect 10226 15076 10232 15088
rect 9806 15048 10232 15076
rect 9806 15045 9818 15048
rect 9760 15039 9818 15045
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18012 15048 18276 15076
rect 18012 15036 18018 15048
rect 11882 15008 11888 15020
rect 9692 14980 11888 15008
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 12158 15008 12164 15020
rect 12115 14980 12164 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12336 15011 12394 15017
rect 12336 14977 12348 15011
rect 12382 15008 12394 15011
rect 13170 15008 13176 15020
rect 12382 14980 13176 15008
rect 12382 14977 12394 14980
rect 12336 14971 12394 14977
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 14636 15011 14694 15017
rect 14636 14977 14648 15011
rect 14682 15008 14694 15011
rect 14918 15008 14924 15020
rect 14682 14980 14924 15008
rect 14682 14977 14694 14980
rect 14636 14971 14694 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 16942 15008 16948 15020
rect 16899 14980 16948 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 17126 15008 17132 15020
rect 17087 14980 17132 15008
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 18138 15008 18144 15020
rect 18099 14980 18144 15008
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18248 15008 18276 15048
rect 18598 15036 18604 15088
rect 18656 15076 18662 15088
rect 20346 15076 20352 15088
rect 18656 15048 19288 15076
rect 18656 15036 18662 15048
rect 19260 15017 19288 15048
rect 19444 15048 20352 15076
rect 19444 15017 19472 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 22094 15076 22100 15088
rect 20456 15048 22100 15076
rect 20456 15017 20484 15048
rect 22094 15036 22100 15048
rect 22152 15036 22158 15088
rect 24317 15023 24345 15116
rect 25590 15104 25596 15116
rect 25648 15104 25654 15156
rect 25958 15104 25964 15156
rect 26016 15144 26022 15156
rect 26421 15147 26479 15153
rect 26421 15144 26433 15147
rect 26016 15116 26433 15144
rect 26016 15104 26022 15116
rect 26421 15113 26433 15116
rect 26467 15113 26479 15147
rect 26421 15107 26479 15113
rect 27706 15104 27712 15156
rect 27764 15144 27770 15156
rect 30650 15144 30656 15156
rect 27764 15116 29684 15144
rect 30611 15116 30656 15144
rect 27764 15104 27770 15116
rect 24946 15076 24952 15088
rect 24412 15048 24952 15076
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18248 14980 18889 15008
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 15008 19671 15011
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 19659 14980 20269 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21266 15008 21272 15020
rect 21223 14980 21272 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 19076 14940 19104 14971
rect 17920 14912 19104 14940
rect 19147 14943 19205 14949
rect 17920 14900 17926 14912
rect 19147 14909 19159 14943
rect 19193 14940 19205 14943
rect 19518 14940 19524 14952
rect 19193 14912 19524 14940
rect 19193 14909 19205 14912
rect 19147 14903 19205 14909
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 20346 14900 20352 14952
rect 20404 14940 20410 14952
rect 20456 14940 20484 14971
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 21818 14968 21824 15020
rect 21876 15008 21882 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21876 14980 22017 15008
rect 21876 14968 21882 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 15008 22523 15011
rect 23474 15008 23480 15020
rect 22511 14980 23480 15008
rect 22511 14977 22523 14980
rect 22465 14971 22523 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 24210 15008 24216 15020
rect 24171 14980 24216 15008
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 24302 15017 24360 15023
rect 24412 15020 24440 15048
rect 24946 15036 24952 15048
rect 25004 15036 25010 15088
rect 25682 15036 25688 15088
rect 25740 15076 25746 15088
rect 27341 15079 27399 15085
rect 27341 15076 27353 15079
rect 25740 15048 27353 15076
rect 25740 15036 25746 15048
rect 27341 15045 27353 15048
rect 27387 15045 27399 15079
rect 27341 15039 27399 15045
rect 27890 15036 27896 15088
rect 27948 15076 27954 15088
rect 29656 15076 29684 15116
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 31297 15147 31355 15153
rect 31297 15144 31309 15147
rect 30760 15116 31309 15144
rect 30760 15076 30788 15116
rect 31297 15113 31309 15116
rect 31343 15113 31355 15147
rect 31297 15107 31355 15113
rect 31202 15076 31208 15088
rect 27948 15048 28212 15076
rect 29656 15048 30788 15076
rect 31163 15048 31208 15076
rect 27948 15036 27954 15048
rect 24302 14983 24314 15017
rect 24348 14983 24360 15017
rect 24302 14977 24360 14983
rect 24397 15014 24455 15020
rect 24397 14980 24409 15014
rect 24443 14980 24455 15014
rect 24397 14974 24455 14980
rect 24581 15011 24639 15017
rect 24581 14977 24593 15011
rect 24627 15008 24639 15011
rect 24670 15008 24676 15020
rect 24627 14980 24676 15008
rect 24627 14977 24639 14980
rect 24581 14971 24639 14977
rect 24670 14968 24676 14980
rect 24728 14968 24734 15020
rect 24854 14968 24860 15020
rect 24912 15008 24918 15020
rect 25314 15017 25320 15020
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24912 14980 25053 15008
rect 24912 14968 24918 14980
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 25297 15011 25320 15017
rect 25297 14977 25309 15011
rect 25297 14971 25320 14977
rect 25314 14968 25320 14971
rect 25372 14968 25378 15020
rect 26970 15008 26976 15020
rect 26931 14980 26976 15008
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 20404 14912 20484 14940
rect 20533 14943 20591 14949
rect 20404 14900 20410 14912
rect 20533 14909 20545 14943
rect 20579 14940 20591 14943
rect 20806 14940 20812 14952
rect 20579 14912 20812 14940
rect 20579 14909 20591 14912
rect 20533 14903 20591 14909
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 22646 14940 22652 14952
rect 20916 14912 22652 14940
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 15436 14844 15761 14872
rect 15436 14832 15442 14844
rect 15749 14841 15761 14844
rect 15795 14872 15807 14875
rect 19426 14872 19432 14884
rect 15795 14844 19432 14872
rect 15795 14841 15807 14844
rect 15749 14835 15807 14841
rect 19426 14832 19432 14844
rect 19484 14872 19490 14884
rect 19886 14872 19892 14884
rect 19484 14844 19892 14872
rect 19484 14832 19490 14844
rect 19886 14832 19892 14844
rect 19944 14832 19950 14884
rect 20070 14872 20076 14884
rect 20031 14844 20076 14872
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 20916 14872 20944 14912
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 23937 14943 23995 14949
rect 22756 14912 23152 14940
rect 20824 14844 20944 14872
rect 10873 14807 10931 14813
rect 10873 14773 10885 14807
rect 10919 14804 10931 14807
rect 11514 14804 11520 14816
rect 10919 14776 11520 14804
rect 10919 14773 10931 14776
rect 10873 14767 10931 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 13136 14776 13461 14804
rect 13136 14764 13142 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 13449 14767 13507 14773
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 18104 14776 18337 14804
rect 18104 14764 18110 14776
rect 18325 14773 18337 14776
rect 18371 14804 18383 14807
rect 20824 14804 20852 14844
rect 21450 14832 21456 14884
rect 21508 14872 21514 14884
rect 22756 14872 22784 14912
rect 21508 14844 22784 14872
rect 22833 14875 22891 14881
rect 21508 14832 21514 14844
rect 22833 14841 22845 14875
rect 22879 14872 22891 14875
rect 23124 14872 23152 14912
rect 23937 14909 23949 14943
rect 23983 14940 23995 14943
rect 24118 14940 24124 14952
rect 23983 14912 24124 14940
rect 23983 14909 23995 14912
rect 23937 14903 23995 14909
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 27172 14940 27200 14971
rect 27982 14968 27988 15020
rect 28040 15008 28046 15020
rect 28184 15017 28212 15048
rect 31202 15036 31208 15048
rect 31260 15036 31266 15088
rect 28077 15011 28135 15017
rect 28077 15008 28089 15011
rect 28040 14980 28089 15008
rect 28040 14968 28046 14980
rect 28077 14977 28089 14980
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28261 15011 28319 15017
rect 28261 14977 28273 15011
rect 28307 14977 28319 15011
rect 28261 14971 28319 14977
rect 26384 14912 27200 14940
rect 28276 14940 28304 14971
rect 28350 14968 28356 15020
rect 28408 15008 28414 15020
rect 28445 15011 28503 15017
rect 28445 15008 28457 15011
rect 28408 14980 28457 15008
rect 28408 14968 28414 14980
rect 28445 14977 28457 14980
rect 28491 14977 28503 15011
rect 29270 15008 29276 15020
rect 29231 14980 29276 15008
rect 28445 14971 28503 14977
rect 29270 14968 29276 14980
rect 29328 14968 29334 15020
rect 29362 14968 29368 15020
rect 29420 15008 29426 15020
rect 29529 15011 29587 15017
rect 29529 15008 29541 15011
rect 29420 14980 29541 15008
rect 29420 14968 29426 14980
rect 29529 14977 29541 14980
rect 29575 14977 29587 15011
rect 29529 14971 29587 14977
rect 29178 14940 29184 14952
rect 28276 14912 29184 14940
rect 26384 14900 26390 14912
rect 29178 14900 29184 14912
rect 29236 14900 29242 14952
rect 25038 14872 25044 14884
rect 22879 14844 23060 14872
rect 23124 14844 25044 14872
rect 22879 14841 22891 14844
rect 22833 14835 22891 14841
rect 20990 14804 20996 14816
rect 18371 14776 20852 14804
rect 20951 14776 20996 14804
rect 18371 14773 18383 14776
rect 18325 14767 18383 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 22925 14807 22983 14813
rect 22925 14804 22937 14807
rect 22704 14776 22937 14804
rect 22704 14764 22710 14776
rect 22925 14773 22937 14776
rect 22971 14773 22983 14807
rect 23032 14804 23060 14844
rect 25038 14832 25044 14844
rect 25096 14832 25102 14884
rect 28810 14872 28816 14884
rect 25976 14844 28816 14872
rect 23198 14804 23204 14816
rect 23032 14776 23204 14804
rect 22925 14767 22983 14773
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 24394 14804 24400 14816
rect 23532 14776 24400 14804
rect 23532 14764 23538 14776
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 25976 14804 26004 14844
rect 28810 14832 28816 14844
rect 28868 14832 28874 14884
rect 24636 14776 26004 14804
rect 27801 14807 27859 14813
rect 24636 14764 24642 14776
rect 27801 14773 27813 14807
rect 27847 14804 27859 14807
rect 29638 14804 29644 14816
rect 27847 14776 29644 14804
rect 27847 14773 27859 14776
rect 27801 14767 27859 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 16114 14600 16120 14612
rect 15703 14572 16120 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 17494 14600 17500 14612
rect 17407 14572 17500 14600
rect 17494 14560 17500 14572
rect 17552 14600 17558 14612
rect 21361 14603 21419 14609
rect 17552 14572 21312 14600
rect 17552 14560 17558 14572
rect 12161 14535 12219 14541
rect 12161 14532 12173 14535
rect 10520 14504 12173 14532
rect 9490 14464 9496 14476
rect 9451 14436 9496 14464
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 9760 14399 9818 14405
rect 9760 14365 9772 14399
rect 9806 14396 9818 14399
rect 10520 14396 10548 14504
rect 12161 14501 12173 14504
rect 12207 14501 12219 14535
rect 12161 14495 12219 14501
rect 17586 14492 17592 14544
rect 17644 14532 17650 14544
rect 19518 14532 19524 14544
rect 17644 14504 19524 14532
rect 17644 14492 17650 14504
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 21284 14532 21312 14572
rect 21361 14569 21373 14603
rect 21407 14600 21419 14603
rect 22278 14600 22284 14612
rect 21407 14572 22284 14600
rect 21407 14569 21419 14572
rect 21361 14563 21419 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 25685 14603 25743 14609
rect 25685 14600 25697 14603
rect 23624 14572 25697 14600
rect 23624 14560 23630 14572
rect 25685 14569 25697 14572
rect 25731 14569 25743 14603
rect 25685 14563 25743 14569
rect 25774 14560 25780 14612
rect 25832 14600 25838 14612
rect 25832 14572 26004 14600
rect 25832 14560 25838 14572
rect 25976 14544 26004 14572
rect 26234 14560 26240 14612
rect 26292 14600 26298 14612
rect 26697 14603 26755 14609
rect 26697 14600 26709 14603
rect 26292 14572 26709 14600
rect 26292 14560 26298 14572
rect 26697 14569 26709 14572
rect 26743 14569 26755 14603
rect 26697 14563 26755 14569
rect 28258 14560 28264 14612
rect 28316 14600 28322 14612
rect 28813 14603 28871 14609
rect 28813 14600 28825 14603
rect 28316 14572 28825 14600
rect 28316 14560 28322 14572
rect 28813 14569 28825 14572
rect 28859 14569 28871 14603
rect 28813 14563 28871 14569
rect 30929 14603 30987 14609
rect 30929 14569 30941 14603
rect 30975 14600 30987 14603
rect 31202 14600 31208 14612
rect 30975 14572 31208 14600
rect 30975 14569 30987 14572
rect 30929 14563 30987 14569
rect 31202 14560 31208 14572
rect 31260 14560 31266 14612
rect 22462 14532 22468 14544
rect 21284 14504 22468 14532
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 25590 14492 25596 14544
rect 25648 14532 25654 14544
rect 25869 14535 25927 14541
rect 25869 14532 25881 14535
rect 25648 14504 25881 14532
rect 25648 14492 25654 14504
rect 25869 14501 25881 14504
rect 25915 14501 25927 14535
rect 25869 14495 25927 14501
rect 25958 14492 25964 14544
rect 26016 14532 26022 14544
rect 26878 14532 26884 14544
rect 26016 14504 26884 14532
rect 26016 14492 26022 14504
rect 26878 14492 26884 14504
rect 26936 14492 26942 14544
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 17862 14464 17868 14476
rect 17184 14436 17868 14464
rect 17184 14424 17190 14436
rect 17862 14424 17868 14436
rect 17920 14464 17926 14476
rect 18325 14467 18383 14473
rect 17920 14436 18184 14464
rect 17920 14424 17926 14436
rect 9806 14368 10548 14396
rect 11701 14399 11759 14405
rect 9806 14365 9818 14368
rect 9760 14359 9818 14365
rect 11701 14365 11713 14399
rect 11747 14396 11759 14399
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 11747 14368 12357 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 14277 14399 14335 14405
rect 12345 14359 12403 14365
rect 12912 14368 14228 14396
rect 12912 14340 12940 14368
rect 11330 14328 11336 14340
rect 11291 14300 11336 14328
rect 11330 14288 11336 14300
rect 11388 14288 11394 14340
rect 11517 14331 11575 14337
rect 11517 14297 11529 14331
rect 11563 14297 11575 14331
rect 12894 14328 12900 14340
rect 12855 14300 12900 14328
rect 11517 14291 11575 14297
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11532 14260 11560 14291
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13113 14331 13171 14337
rect 13113 14297 13125 14331
rect 13159 14328 13171 14331
rect 13446 14328 13452 14340
rect 13159 14300 13452 14328
rect 13159 14297 13171 14300
rect 13113 14291 13171 14297
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 13262 14260 13268 14272
rect 10919 14232 11560 14260
rect 13223 14232 13268 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 14200 14260 14228 14368
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 14366 14396 14372 14408
rect 14323 14368 14372 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 14366 14356 14372 14368
rect 14424 14396 14430 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 14424 14368 16129 14396
rect 14424 14356 14430 14368
rect 16117 14365 16129 14368
rect 16163 14396 16175 14399
rect 16206 14396 16212 14408
rect 16163 14368 16212 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 17954 14396 17960 14408
rect 17915 14368 17960 14396
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18156 14405 18184 14436
rect 18325 14433 18337 14467
rect 18371 14464 18383 14467
rect 18598 14464 18604 14476
rect 18371 14436 18604 14464
rect 18371 14433 18383 14436
rect 18325 14427 18383 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19978 14464 19984 14476
rect 19939 14436 19984 14464
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 21008 14436 27476 14464
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18414 14396 18420 14408
rect 18279 14368 18420 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18690 14396 18696 14408
rect 18555 14368 18696 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 20622 14396 20628 14408
rect 19484 14368 20628 14396
rect 19484 14356 19490 14368
rect 20622 14356 20628 14368
rect 20680 14396 20686 14408
rect 21008 14396 21036 14436
rect 20680 14368 21036 14396
rect 20680 14356 20686 14368
rect 21542 14356 21548 14408
rect 21600 14396 21606 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21600 14368 21833 14396
rect 21600 14356 21606 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14396 22063 14399
rect 22094 14396 22100 14408
rect 22051 14368 22100 14396
rect 22051 14365 22063 14368
rect 22005 14359 22063 14365
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22646 14396 22652 14408
rect 22244 14368 22324 14396
rect 22607 14368 22652 14396
rect 22244 14356 22250 14368
rect 14544 14331 14602 14337
rect 14544 14297 14556 14331
rect 14590 14328 14602 14331
rect 15286 14328 15292 14340
rect 14590 14300 15292 14328
rect 14590 14297 14602 14300
rect 14544 14291 14602 14297
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 16384 14331 16442 14337
rect 16384 14297 16396 14331
rect 16430 14328 16442 14331
rect 16666 14328 16672 14340
rect 16430 14300 16672 14328
rect 16430 14297 16442 14300
rect 16384 14291 16442 14297
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 19337 14331 19395 14337
rect 19337 14328 19349 14331
rect 18156 14300 19349 14328
rect 18156 14272 18184 14300
rect 19337 14297 19349 14300
rect 19383 14297 19395 14331
rect 19337 14291 19395 14297
rect 20248 14331 20306 14337
rect 20248 14297 20260 14331
rect 20294 14328 20306 14331
rect 20898 14328 20904 14340
rect 20294 14300 20904 14328
rect 20294 14297 20306 14300
rect 20248 14291 20306 14297
rect 20898 14288 20904 14300
rect 20956 14288 20962 14340
rect 15654 14260 15660 14272
rect 14200 14232 15660 14260
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 18138 14220 18144 14272
rect 18196 14220 18202 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18472 14232 18705 14260
rect 18472 14220 18478 14232
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 19429 14263 19487 14269
rect 19429 14229 19441 14263
rect 19475 14260 19487 14263
rect 22002 14260 22008 14272
rect 19475 14232 22008 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 22186 14260 22192 14272
rect 22147 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22296 14260 22324 14368
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 22796 14368 22841 14396
rect 22796 14356 22802 14368
rect 23106 14356 23112 14408
rect 23164 14405 23170 14408
rect 23164 14396 23172 14405
rect 24394 14396 24400 14408
rect 23164 14368 23209 14396
rect 24355 14368 24400 14396
rect 23164 14359 23172 14368
rect 23164 14356 23170 14359
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 24490 14399 24548 14405
rect 24490 14365 24502 14399
rect 24536 14365 24548 14399
rect 24670 14396 24676 14408
rect 24631 14368 24676 14396
rect 24490 14359 24548 14365
rect 22922 14328 22928 14340
rect 22883 14300 22928 14328
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 23017 14331 23075 14337
rect 23017 14297 23029 14331
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 23032 14260 23060 14291
rect 23842 14288 23848 14340
rect 23900 14328 23906 14340
rect 24504 14328 24532 14359
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 24862 14399 24920 14405
rect 24862 14365 24874 14399
rect 24908 14396 24920 14399
rect 24908 14368 24992 14396
rect 24908 14365 24920 14368
rect 24862 14359 24920 14365
rect 23900 14300 24532 14328
rect 23900 14288 23906 14300
rect 24762 14288 24768 14340
rect 24820 14328 24826 14340
rect 24964 14328 24992 14368
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 27448 14405 27476 14436
rect 27798 14424 27804 14476
rect 27856 14464 27862 14476
rect 28534 14464 28540 14476
rect 27856 14436 28540 14464
rect 27856 14424 27862 14436
rect 28534 14424 28540 14436
rect 28592 14464 28598 14476
rect 28592 14436 28764 14464
rect 28592 14424 28598 14436
rect 27433 14399 27491 14405
rect 25096 14368 25544 14396
rect 25096 14356 25102 14368
rect 25516 14337 25544 14368
rect 27433 14365 27445 14399
rect 27479 14365 27491 14399
rect 27614 14396 27620 14408
rect 27575 14368 27620 14396
rect 27433 14359 27491 14365
rect 27614 14356 27620 14368
rect 27672 14396 27678 14408
rect 28736 14405 28764 14436
rect 29270 14424 29276 14476
rect 29328 14464 29334 14476
rect 29549 14467 29607 14473
rect 29549 14464 29561 14467
rect 29328 14436 29561 14464
rect 29328 14424 29334 14436
rect 29549 14433 29561 14436
rect 29595 14433 29607 14467
rect 29549 14427 29607 14433
rect 28261 14399 28319 14405
rect 27672 14368 28212 14396
rect 27672 14356 27678 14368
rect 25501 14331 25559 14337
rect 24820 14300 24865 14328
rect 24964 14300 25176 14328
rect 24820 14288 24826 14300
rect 23290 14260 23296 14272
rect 22296 14232 23060 14260
rect 23251 14232 23296 14260
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 25041 14263 25099 14269
rect 25041 14260 25053 14263
rect 24912 14232 25053 14260
rect 24912 14220 24918 14232
rect 25041 14229 25053 14232
rect 25087 14229 25099 14263
rect 25148 14260 25176 14300
rect 25501 14297 25513 14331
rect 25547 14297 25559 14331
rect 26513 14331 26571 14337
rect 25501 14291 25559 14297
rect 25792 14300 26004 14328
rect 25682 14260 25688 14272
rect 25740 14269 25746 14272
rect 25740 14263 25759 14269
rect 25148 14232 25688 14260
rect 25041 14223 25099 14229
rect 25682 14220 25688 14232
rect 25747 14260 25759 14263
rect 25792 14260 25820 14300
rect 25747 14232 25820 14260
rect 25976 14260 26004 14300
rect 26513 14297 26525 14331
rect 26559 14328 26571 14331
rect 27706 14328 27712 14340
rect 26559 14300 27712 14328
rect 26559 14297 26571 14300
rect 26513 14291 26571 14297
rect 27706 14288 27712 14300
rect 27764 14288 27770 14340
rect 26713 14263 26771 14269
rect 26713 14260 26725 14263
rect 25976 14232 26725 14260
rect 25747 14229 25759 14232
rect 25740 14223 25759 14229
rect 26713 14229 26725 14232
rect 26759 14229 26771 14263
rect 26878 14260 26884 14272
rect 26839 14232 26884 14260
rect 26713 14223 26771 14229
rect 25740 14220 25746 14223
rect 26878 14220 26884 14232
rect 26936 14220 26942 14272
rect 27430 14220 27436 14272
rect 27488 14260 27494 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27488 14232 28089 14260
rect 27488 14220 27494 14232
rect 28077 14229 28089 14232
rect 28123 14229 28135 14263
rect 28184 14260 28212 14368
rect 28261 14365 28273 14399
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28902 14396 28908 14408
rect 28863 14368 28908 14396
rect 28721 14359 28779 14365
rect 28276 14328 28304 14359
rect 28902 14356 28908 14368
rect 28960 14356 28966 14408
rect 29638 14356 29644 14408
rect 29696 14396 29702 14408
rect 29805 14399 29863 14405
rect 29805 14396 29817 14399
rect 29696 14368 29817 14396
rect 29696 14356 29702 14368
rect 29805 14365 29817 14368
rect 29851 14365 29863 14399
rect 29805 14359 29863 14365
rect 29086 14328 29092 14340
rect 28276 14300 29092 14328
rect 29086 14288 29092 14300
rect 29144 14288 29150 14340
rect 28350 14260 28356 14272
rect 28184 14232 28356 14260
rect 28077 14223 28135 14229
rect 28350 14220 28356 14232
rect 28408 14220 28414 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 8849 14059 8907 14065
rect 8849 14025 8861 14059
rect 8895 14056 8907 14059
rect 9766 14056 9772 14068
rect 8895 14028 9772 14056
rect 8895 14025 8907 14028
rect 8849 14019 8907 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10873 14059 10931 14065
rect 10873 14025 10885 14059
rect 10919 14056 10931 14059
rect 10919 14028 11744 14056
rect 10919 14025 10931 14028
rect 10873 14019 10931 14025
rect 10502 13988 10508 14000
rect 9048 13960 10508 13988
rect 9048 13929 9076 13960
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 11716 13997 11744 14028
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 11940 14028 12725 14056
rect 11940 14016 11946 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 12713 14019 12771 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 14918 14056 14924 14068
rect 14879 14028 14924 14056
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 16666 14056 16672 14068
rect 16627 14028 16672 14056
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 18230 14056 18236 14068
rect 17788 14028 18236 14056
rect 11701 13991 11759 13997
rect 11701 13957 11713 13991
rect 11747 13957 11759 13991
rect 11701 13951 11759 13957
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 12529 13991 12587 13997
rect 12529 13988 12541 13991
rect 11848 13960 12541 13988
rect 11848 13948 11854 13960
rect 12529 13957 12541 13960
rect 12575 13957 12587 13991
rect 12529 13951 12587 13957
rect 16117 13991 16175 13997
rect 16117 13957 16129 13991
rect 16163 13988 16175 13991
rect 16390 13988 16396 14000
rect 16163 13960 16396 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17788 13988 17816 14028
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 18340 14028 19472 14056
rect 16684 13960 17816 13988
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9760 13923 9818 13929
rect 9760 13889 9772 13923
rect 9806 13920 9818 13923
rect 10226 13920 10232 13932
rect 9806 13892 10232 13920
rect 9806 13889 9818 13892
rect 9760 13883 9818 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11388 13892 11529 13920
rect 11388 13880 11394 13892
rect 11517 13889 11529 13892
rect 11563 13920 11575 13923
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 11563 13892 12357 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13320 13892 13369 13920
rect 13320 13880 13326 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 14550 13920 14556 13932
rect 14507 13892 14556 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15194 13920 15200 13932
rect 15151 13892 15200 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15933 13923 15991 13929
rect 15335 13892 15516 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 9490 13852 9496 13864
rect 9451 13824 9496 13852
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 15378 13852 15384 13864
rect 15339 13824 15384 13852
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15488 13852 15516 13892
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16684 13920 16712 13960
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18340 13988 18368 14028
rect 18690 13988 18696 14000
rect 17920 13960 18368 13988
rect 17920 13948 17926 13960
rect 16850 13920 16856 13932
rect 15979 13892 16712 13920
rect 16811 13892 16856 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17494 13920 17500 13932
rect 17175 13892 17500 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 17644 13892 18061 13920
rect 17644 13880 17650 13892
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13920 18291 13923
rect 18340 13920 18368 13960
rect 18432 13960 18696 13988
rect 18432 13929 18460 13960
rect 18690 13948 18696 13960
rect 18748 13988 18754 14000
rect 18748 13960 19380 13988
rect 18748 13948 18754 13960
rect 18279 13892 18368 13920
rect 18417 13923 18475 13929
rect 18279 13889 18291 13892
rect 18233 13883 18291 13889
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13920 18659 13923
rect 18966 13920 18972 13932
rect 18647 13892 18972 13920
rect 18647 13889 18659 13892
rect 18601 13883 18659 13889
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 15746 13852 15752 13864
rect 15488 13824 15752 13852
rect 15746 13812 15752 13824
rect 15804 13852 15810 13864
rect 17037 13855 17095 13861
rect 17037 13852 17049 13855
rect 15804 13824 17049 13852
rect 15804 13812 15810 13824
rect 17037 13821 17049 13824
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 18012 13824 18337 13852
rect 18012 13812 18018 13824
rect 18325 13821 18337 13824
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 19058 13784 19064 13796
rect 17184 13756 19064 13784
rect 17184 13744 17190 13756
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 19260 13784 19288 13883
rect 19352 13852 19380 13960
rect 19444 13935 19472 14028
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20622 14056 20628 14068
rect 20404 14028 20628 14056
rect 20404 14016 20410 14028
rect 20622 14016 20628 14028
rect 20680 14056 20686 14068
rect 20680 14028 20760 14056
rect 20680 14016 20686 14028
rect 19429 13929 19487 13935
rect 19429 13895 19441 13929
rect 19475 13895 19487 13929
rect 19429 13889 19487 13895
rect 19518 13880 19524 13932
rect 19576 13920 19582 13932
rect 19797 13923 19855 13929
rect 19576 13892 19621 13920
rect 19576 13880 19582 13892
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 20162 13920 20168 13932
rect 19843 13892 20168 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20404 13892 20637 13920
rect 20404 13880 20410 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20732 13920 20760 14028
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 22649 14059 22707 14065
rect 22649 14056 22661 14059
rect 20864 14028 22661 14056
rect 20864 14016 20870 14028
rect 22649 14025 22661 14028
rect 22695 14025 22707 14059
rect 22649 14019 22707 14025
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 24578 14056 24584 14068
rect 24360 14028 24584 14056
rect 24360 14016 24366 14028
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 25148 14028 28549 14056
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22244 13960 24808 13988
rect 22244 13948 22250 13960
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20732 13892 20821 13920
rect 20625 13883 20683 13889
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21784 13892 21833 13920
rect 21784 13880 21790 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 22002 13920 22008 13932
rect 21963 13892 22008 13920
rect 21821 13883 21879 13889
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 22830 13920 22836 13932
rect 22791 13892 22836 13920
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 24780 13929 24808 13960
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 24854 13880 24860 13932
rect 24912 13920 24918 13932
rect 25148 13929 25176 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 29178 14016 29184 14068
rect 29236 14056 29242 14068
rect 29733 14059 29791 14065
rect 29733 14056 29745 14059
rect 29236 14028 29745 14056
rect 29236 14016 29242 14028
rect 29733 14025 29745 14028
rect 29779 14025 29791 14059
rect 29733 14019 29791 14025
rect 26050 13988 26056 14000
rect 26011 13960 26056 13988
rect 26050 13948 26056 13960
rect 26108 13948 26114 14000
rect 26253 13991 26311 13997
rect 26253 13988 26265 13991
rect 26160 13960 26265 13988
rect 25133 13923 25191 13929
rect 24912 13892 24957 13920
rect 24912 13880 24918 13892
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 26160 13920 26188 13960
rect 26253 13957 26265 13960
rect 26299 13957 26311 13991
rect 28626 13988 28632 14000
rect 26253 13951 26311 13957
rect 27172 13960 28632 13988
rect 27172 13929 27200 13960
rect 28626 13948 28632 13960
rect 28684 13948 28690 14000
rect 28718 13948 28724 14000
rect 28776 13988 28782 14000
rect 28776 13960 29868 13988
rect 28776 13948 28782 13960
rect 27430 13929 27436 13932
rect 25133 13883 25191 13889
rect 25700 13892 26188 13920
rect 27157 13923 27215 13929
rect 25700 13864 25728 13892
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27424 13920 27436 13929
rect 27391 13892 27436 13920
rect 27157 13883 27215 13889
rect 27424 13883 27436 13892
rect 27430 13880 27436 13883
rect 27488 13880 27494 13932
rect 29178 13920 29184 13932
rect 29139 13892 29184 13920
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 29840 13929 29868 13960
rect 29641 13923 29699 13929
rect 29641 13889 29653 13923
rect 29687 13889 29699 13923
rect 29641 13883 29699 13889
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13889 29883 13923
rect 29825 13883 29883 13889
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19352 13824 19625 13852
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 20530 13812 20536 13864
rect 20588 13852 20594 13864
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20588 13824 20913 13852
rect 20588 13812 20594 13824
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 22189 13855 22247 13861
rect 22189 13821 22201 13855
rect 22235 13852 22247 13855
rect 22646 13852 22652 13864
rect 22235 13824 22652 13852
rect 22235 13821 22247 13824
rect 22189 13815 22247 13821
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 22922 13852 22928 13864
rect 22796 13824 22928 13852
rect 22796 13812 22802 13824
rect 22922 13812 22928 13824
rect 22980 13852 22986 13864
rect 23293 13855 23351 13861
rect 23293 13852 23305 13855
rect 22980 13824 23305 13852
rect 22980 13812 22986 13824
rect 23293 13821 23305 13824
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 23569 13855 23627 13861
rect 23569 13821 23581 13855
rect 23615 13852 23627 13855
rect 25682 13852 25688 13864
rect 23615 13824 25688 13852
rect 23615 13821 23627 13824
rect 23569 13815 23627 13821
rect 24872 13796 24900 13824
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 28534 13812 28540 13864
rect 28592 13852 28598 13864
rect 29656 13852 29684 13883
rect 28592 13824 29684 13852
rect 28592 13812 28598 13824
rect 19260 13756 19656 13784
rect 19628 13728 19656 13756
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 20441 13787 20499 13793
rect 20441 13784 20453 13787
rect 20128 13756 20453 13784
rect 20128 13744 20134 13756
rect 20441 13753 20453 13756
rect 20487 13753 20499 13787
rect 20441 13747 20499 13753
rect 22462 13744 22468 13796
rect 22520 13784 22526 13796
rect 23014 13784 23020 13796
rect 22520 13756 23020 13784
rect 22520 13744 22526 13756
rect 23014 13744 23020 13756
rect 23072 13744 23078 13796
rect 23198 13744 23204 13796
rect 23256 13784 23262 13796
rect 24670 13784 24676 13796
rect 23256 13756 24676 13784
rect 23256 13744 23262 13756
rect 24670 13744 24676 13756
rect 24728 13744 24734 13796
rect 24854 13744 24860 13796
rect 24912 13744 24918 13796
rect 25041 13787 25099 13793
rect 25041 13753 25053 13787
rect 25087 13784 25099 13787
rect 25130 13784 25136 13796
rect 25087 13756 25136 13784
rect 25087 13753 25099 13756
rect 25041 13747 25099 13753
rect 25130 13744 25136 13756
rect 25188 13744 25194 13796
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11112 13688 11897 13716
rect 11112 13676 11118 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 14274 13716 14280 13728
rect 14235 13688 14280 13716
rect 11885 13679 11943 13685
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 17678 13676 17684 13728
rect 17736 13716 17742 13728
rect 17862 13716 17868 13728
rect 17736 13688 17868 13716
rect 17736 13676 17742 13688
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 18785 13719 18843 13725
rect 18785 13716 18797 13719
rect 18748 13688 18797 13716
rect 18748 13676 18754 13688
rect 18785 13685 18797 13688
rect 18831 13685 18843 13719
rect 18785 13679 18843 13685
rect 18874 13676 18880 13728
rect 18932 13716 18938 13728
rect 19242 13716 19248 13728
rect 18932 13688 19248 13716
rect 18932 13676 18938 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19610 13676 19616 13728
rect 19668 13676 19674 13728
rect 19981 13719 20039 13725
rect 19981 13685 19993 13719
rect 20027 13716 20039 13719
rect 20254 13716 20260 13728
rect 20027 13688 20260 13716
rect 20027 13685 20039 13688
rect 19981 13679 20039 13685
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 23382 13676 23388 13728
rect 23440 13716 23446 13728
rect 25222 13716 25228 13728
rect 23440 13688 25228 13716
rect 23440 13676 23446 13688
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 25314 13676 25320 13728
rect 25372 13716 25378 13728
rect 26234 13716 26240 13728
rect 25372 13688 26240 13716
rect 25372 13676 25378 13688
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 26421 13719 26479 13725
rect 26421 13685 26433 13719
rect 26467 13716 26479 13719
rect 26970 13716 26976 13728
rect 26467 13688 26976 13716
rect 26467 13685 26479 13688
rect 26421 13679 26479 13685
rect 26970 13676 26976 13688
rect 27028 13676 27034 13728
rect 28994 13716 29000 13728
rect 28955 13688 29000 13716
rect 28994 13676 29000 13688
rect 29052 13676 29058 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 10962 13512 10968 13524
rect 10919 13484 10968 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 19978 13512 19984 13524
rect 19720 13484 19984 13512
rect 13354 13444 13360 13456
rect 13315 13416 13360 13444
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 17218 13444 17224 13456
rect 17179 13416 17224 13444
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 17678 13404 17684 13456
rect 17736 13444 17742 13456
rect 17736 13416 19555 13444
rect 17736 13404 17742 13416
rect 19426 13376 19432 13388
rect 13188 13348 19432 13376
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9490 13308 9496 13320
rect 9088 13280 9496 13308
rect 9088 13268 9094 13280
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9766 13317 9772 13320
rect 9760 13308 9772 13317
rect 9727 13280 9772 13308
rect 9760 13271 9772 13280
rect 9766 13268 9772 13271
rect 9824 13268 9830 13320
rect 11514 13308 11520 13320
rect 11475 13280 11520 13308
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 13188 13317 13216 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 12032 13280 12265 13308
rect 12032 13268 12038 13280
rect 12253 13277 12265 13280
rect 12299 13308 12311 13311
rect 13173 13311 13231 13317
rect 12299 13280 13124 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 11330 13240 11336 13252
rect 11291 13212 11336 13240
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 12986 13240 12992 13252
rect 12483 13212 12992 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 13096 13240 13124 13280
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 13998 13308 14004 13320
rect 13688 13280 14004 13308
rect 13688 13268 13694 13280
rect 13998 13268 14004 13280
rect 14056 13308 14062 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 14056 13280 14105 13308
rect 14056 13268 14062 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14918 13308 14924 13320
rect 14879 13280 14924 13308
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 13096 13212 14197 13240
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 15580 13240 15608 13271
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15896 13280 16221 13308
rect 15896 13268 15902 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13308 17095 13311
rect 18138 13308 18144 13320
rect 17083 13280 18144 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18414 13308 18420 13320
rect 18375 13280 18420 13308
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13308 18751 13311
rect 19334 13308 19340 13320
rect 18739 13280 19340 13308
rect 18739 13277 18751 13280
rect 18693 13271 18751 13277
rect 14185 13203 14243 13209
rect 14292 13212 15608 13240
rect 18616 13240 18644 13271
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19527 13308 19555 13416
rect 19720 13385 19748 13484
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 21085 13515 21143 13521
rect 21085 13512 21097 13515
rect 21048 13484 21097 13512
rect 21048 13472 21054 13484
rect 21085 13481 21097 13484
rect 21131 13481 21143 13515
rect 21085 13475 21143 13481
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 24486 13512 24492 13524
rect 23164 13484 23336 13512
rect 23164 13472 23170 13484
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 22152 13348 22600 13376
rect 22152 13336 22158 13348
rect 21266 13308 21272 13320
rect 19527 13280 21272 13308
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 22462 13308 22468 13320
rect 22423 13280 22468 13308
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 22572 13308 22600 13348
rect 22922 13336 22928 13388
rect 22980 13376 22986 13388
rect 23308 13385 23336 13484
rect 23584 13484 24492 13512
rect 23201 13379 23259 13385
rect 23201 13376 23213 13379
rect 22980 13348 23213 13376
rect 22980 13336 22986 13348
rect 23201 13345 23213 13348
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 23584 13317 23612 13484
rect 24486 13472 24492 13484
rect 24544 13512 24550 13524
rect 25685 13515 25743 13521
rect 25685 13512 25697 13515
rect 24544 13484 25697 13512
rect 24544 13472 24550 13484
rect 25685 13481 25697 13484
rect 25731 13481 25743 13515
rect 25685 13475 25743 13481
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 28169 13515 28227 13521
rect 26476 13484 27016 13512
rect 26476 13472 26482 13484
rect 24210 13404 24216 13456
rect 24268 13444 24274 13456
rect 24268 13416 24717 13444
rect 24268 13404 24274 13416
rect 24118 13336 24124 13388
rect 24176 13376 24182 13388
rect 24689 13376 24717 13416
rect 24762 13404 24768 13456
rect 24820 13444 24826 13456
rect 25041 13447 25099 13453
rect 25041 13444 25053 13447
rect 24820 13416 25053 13444
rect 24820 13404 24826 13416
rect 25041 13413 25053 13416
rect 25087 13413 25099 13447
rect 25041 13407 25099 13413
rect 26878 13404 26884 13456
rect 26936 13404 26942 13456
rect 24176 13348 24533 13376
rect 24689 13348 24808 13376
rect 24176 13336 24182 13348
rect 23109 13311 23167 13317
rect 23109 13308 23121 13311
rect 22572 13280 23121 13308
rect 23109 13277 23121 13280
rect 23155 13277 23167 13311
rect 23109 13271 23167 13277
rect 23385 13311 23443 13317
rect 23385 13277 23397 13311
rect 23431 13277 23443 13311
rect 23385 13271 23443 13277
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 23569 13271 23627 13277
rect 19972 13243 20030 13249
rect 18616 13212 18736 13240
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14292 13172 14320 13212
rect 14734 13172 14740 13184
rect 13872 13144 14320 13172
rect 14695 13144 14740 13172
rect 13872 13132 13878 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 15378 13172 15384 13184
rect 15339 13144 15384 13172
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 16025 13175 16083 13181
rect 16025 13172 16037 13175
rect 15988 13144 16037 13172
rect 15988 13132 15994 13144
rect 16025 13141 16037 13144
rect 16071 13141 16083 13175
rect 18230 13172 18236 13184
rect 18191 13144 18236 13172
rect 16025 13135 16083 13141
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 18708 13172 18736 13212
rect 19972 13209 19984 13243
rect 20018 13240 20030 13243
rect 20070 13240 20076 13252
rect 20018 13212 20076 13240
rect 20018 13209 20030 13212
rect 19972 13203 20030 13209
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 22005 13243 22063 13249
rect 22005 13209 22017 13243
rect 22051 13240 22063 13243
rect 23400 13240 23428 13271
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24505 13317 24533 13348
rect 24490 13311 24548 13317
rect 24490 13277 24502 13311
rect 24536 13277 24548 13311
rect 24670 13308 24676 13320
rect 24631 13280 24676 13308
rect 24490 13271 24548 13277
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 24780 13317 24808 13348
rect 24946 13336 24952 13388
rect 25004 13376 25010 13388
rect 26896 13376 26924 13404
rect 25004 13348 25544 13376
rect 25004 13336 25010 13348
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24854 13268 24860 13320
rect 24912 13317 24918 13320
rect 25516 13317 25544 13348
rect 26712 13348 26924 13376
rect 24912 13308 24920 13317
rect 25501 13311 25559 13317
rect 24912 13280 24957 13308
rect 24912 13271 24920 13280
rect 25501 13277 25513 13311
rect 25547 13308 25559 13311
rect 25590 13308 25596 13320
rect 25547 13280 25596 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 24912 13268 24918 13271
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 26712 13317 26740 13348
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 26845 13311 26903 13317
rect 26845 13277 26857 13311
rect 26891 13308 26903 13311
rect 26988 13308 27016 13484
rect 28169 13481 28181 13515
rect 28215 13512 28227 13515
rect 29178 13512 29184 13524
rect 28215 13484 29184 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 29178 13472 29184 13484
rect 29236 13472 29242 13524
rect 28997 13447 29055 13453
rect 28997 13413 29009 13447
rect 29043 13444 29055 13447
rect 29086 13444 29092 13456
rect 29043 13416 29092 13444
rect 29043 13413 29055 13416
rect 28997 13407 29055 13413
rect 29086 13404 29092 13416
rect 29144 13404 29150 13456
rect 27246 13317 27252 13320
rect 26891 13280 27016 13308
rect 27203 13311 27252 13317
rect 26891 13277 26903 13280
rect 26845 13271 26903 13277
rect 27203 13277 27215 13311
rect 27249 13277 27252 13311
rect 27203 13271 27252 13277
rect 27246 13268 27252 13271
rect 27304 13268 27310 13320
rect 28629 13311 28687 13317
rect 28629 13308 28641 13311
rect 27816 13280 28641 13308
rect 22051 13212 23428 13240
rect 22051 13209 22063 13212
rect 22005 13203 22063 13209
rect 26418 13200 26424 13252
rect 26476 13240 26482 13252
rect 26973 13243 27031 13249
rect 26973 13240 26985 13243
rect 26476 13212 26985 13240
rect 26476 13200 26482 13212
rect 26973 13209 26985 13212
rect 27019 13209 27031 13243
rect 26973 13203 27031 13209
rect 27065 13243 27123 13249
rect 27065 13209 27077 13243
rect 27111 13240 27123 13243
rect 27111 13212 27660 13240
rect 27111 13209 27123 13212
rect 27065 13203 27123 13209
rect 20622 13172 20628 13184
rect 18708 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 22373 13175 22431 13181
rect 22373 13141 22385 13175
rect 22419 13172 22431 13175
rect 22462 13172 22468 13184
rect 22419 13144 22468 13172
rect 22419 13141 22431 13144
rect 22373 13135 22431 13141
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 22925 13175 22983 13181
rect 22925 13141 22937 13175
rect 22971 13172 22983 13175
rect 23014 13172 23020 13184
rect 22971 13144 23020 13172
rect 22971 13141 22983 13144
rect 22925 13135 22983 13141
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 27341 13175 27399 13181
rect 27341 13141 27353 13175
rect 27387 13172 27399 13175
rect 27522 13172 27528 13184
rect 27387 13144 27528 13172
rect 27387 13141 27399 13144
rect 27341 13135 27399 13141
rect 27522 13132 27528 13144
rect 27580 13132 27586 13184
rect 27632 13172 27660 13212
rect 27706 13200 27712 13252
rect 27764 13240 27770 13252
rect 27816 13249 27844 13280
rect 28629 13277 28641 13280
rect 28675 13277 28687 13311
rect 28810 13308 28816 13320
rect 28771 13280 28816 13308
rect 28629 13271 28687 13277
rect 28810 13268 28816 13280
rect 28868 13268 28874 13320
rect 27801 13243 27859 13249
rect 27801 13240 27813 13243
rect 27764 13212 27813 13240
rect 27764 13200 27770 13212
rect 27801 13209 27813 13212
rect 27847 13209 27859 13243
rect 27801 13203 27859 13209
rect 27890 13200 27896 13252
rect 27948 13240 27954 13252
rect 27985 13243 28043 13249
rect 27985 13240 27997 13243
rect 27948 13212 27997 13240
rect 27948 13200 27954 13212
rect 27985 13209 27997 13212
rect 28031 13209 28043 13243
rect 27985 13203 28043 13209
rect 28902 13172 28908 13184
rect 27632 13144 28908 13172
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 10226 12968 10232 12980
rect 10187 12940 10232 12968
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 12986 12968 12992 12980
rect 12947 12940 12992 12968
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14458 12968 14464 12980
rect 14056 12940 14464 12968
rect 14056 12928 14062 12940
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 14826 12968 14832 12980
rect 14787 12940 14832 12968
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 20070 12968 20076 12980
rect 17092 12940 18552 12968
rect 20031 12940 20076 12968
rect 17092 12928 17098 12940
rect 11876 12903 11934 12909
rect 11876 12869 11888 12903
rect 11922 12900 11934 12903
rect 12434 12900 12440 12912
rect 11922 12872 12440 12900
rect 11922 12869 11934 12872
rect 11876 12863 11934 12869
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 13716 12903 13774 12909
rect 13716 12869 13728 12903
rect 13762 12900 13774 12903
rect 14734 12900 14740 12912
rect 13762 12872 14740 12900
rect 13762 12869 13774 12872
rect 13716 12863 13774 12869
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 16942 12860 16948 12912
rect 17000 12900 17006 12912
rect 17000 12872 18184 12900
rect 17000 12860 17006 12872
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 11054 12832 11060 12844
rect 10459 12804 11060 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 9784 12764 9812 12795
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 12216 12804 13461 12832
rect 12216 12792 12222 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 15470 12832 15476 12844
rect 15431 12804 15476 12832
rect 13449 12795 13507 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 15746 12792 15752 12844
rect 15804 12832 15810 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15804 12804 16129 12832
rect 15804 12792 15810 12804
rect 16117 12801 16129 12804
rect 16163 12801 16175 12835
rect 16850 12832 16856 12844
rect 16811 12804 16856 12832
rect 16117 12795 16175 12801
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17681 12835 17739 12841
rect 17681 12832 17693 12835
rect 17083 12804 17693 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17681 12801 17693 12804
rect 17727 12801 17739 12835
rect 18156 12832 18184 12872
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 18386 12903 18444 12909
rect 18386 12900 18398 12903
rect 18288 12872 18398 12900
rect 18288 12860 18294 12872
rect 18386 12869 18398 12872
rect 18432 12869 18444 12903
rect 18524 12900 18552 12940
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 21140 12940 21864 12968
rect 21140 12928 21146 12940
rect 18524 12872 21772 12900
rect 18386 12863 18444 12869
rect 19426 12832 19432 12844
rect 18156 12804 19432 12832
rect 17681 12795 17739 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20441 12835 20499 12841
rect 20441 12801 20453 12835
rect 20487 12832 20499 12835
rect 20622 12832 20628 12844
rect 20487 12804 20628 12832
rect 20487 12801 20499 12804
rect 20441 12795 20499 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21266 12832 21272 12844
rect 21227 12804 21272 12832
rect 21085 12795 21143 12801
rect 11422 12764 11428 12776
rect 9784 12736 11428 12764
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11606 12764 11612 12776
rect 11567 12736 11612 12764
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 18046 12764 18052 12776
rect 16715 12736 18052 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18141 12767 18199 12773
rect 18141 12733 18153 12767
rect 18187 12733 18199 12767
rect 18141 12727 18199 12733
rect 20533 12767 20591 12773
rect 20533 12733 20545 12767
rect 20579 12764 20591 12767
rect 20990 12764 20996 12776
rect 20579 12736 20996 12764
rect 20579 12733 20591 12736
rect 20533 12727 20591 12733
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10962 12696 10968 12708
rect 9631 12668 10968 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 15933 12699 15991 12705
rect 15933 12696 15945 12699
rect 14384 12668 15945 12696
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 14384 12628 14412 12668
rect 15933 12665 15945 12668
rect 15979 12665 15991 12699
rect 15933 12659 15991 12665
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 18156 12696 18184 12727
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21100 12764 21128 12795
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 21634 12764 21640 12776
rect 21100 12736 21640 12764
rect 21634 12724 21640 12736
rect 21692 12724 21698 12776
rect 21744 12764 21772 12872
rect 21836 12841 21864 12940
rect 22462 12928 22468 12980
rect 22520 12968 22526 12980
rect 22520 12940 22968 12968
rect 22520 12928 22526 12940
rect 22830 12900 22836 12912
rect 21928 12872 22836 12900
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 21928 12764 21956 12872
rect 22830 12860 22836 12872
rect 22888 12860 22894 12912
rect 22940 12900 22968 12940
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 23532 12940 25237 12968
rect 23532 12928 23538 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 30009 12971 30067 12977
rect 30009 12968 30021 12971
rect 25225 12931 25283 12937
rect 27356 12940 30021 12968
rect 23750 12900 23756 12912
rect 22940 12872 23756 12900
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 24949 12903 25007 12909
rect 24949 12869 24961 12903
rect 24995 12900 25007 12903
rect 25498 12900 25504 12912
rect 24995 12872 25504 12900
rect 24995 12869 25007 12872
rect 24949 12863 25007 12869
rect 25498 12860 25504 12872
rect 25556 12860 25562 12912
rect 25682 12900 25688 12912
rect 25643 12872 25688 12900
rect 25682 12860 25688 12872
rect 25740 12860 25746 12912
rect 25885 12903 25943 12909
rect 25885 12900 25897 12903
rect 25792 12872 25897 12900
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 23014 12841 23020 12844
rect 23008 12832 23020 12841
rect 22060 12804 22105 12832
rect 22975 12804 23020 12832
rect 22060 12792 22066 12804
rect 23008 12795 23020 12804
rect 23014 12792 23020 12795
rect 23072 12792 23078 12844
rect 21744 12736 21956 12764
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22520 12736 22753 12764
rect 22520 12724 22526 12736
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 23768 12764 23796 12860
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24452 12804 24593 12832
rect 24452 12792 24458 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 24674 12835 24732 12841
rect 24674 12801 24686 12835
rect 24720 12801 24732 12835
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 24674 12795 24732 12801
rect 24771 12804 24869 12832
rect 24688 12764 24716 12795
rect 23768 12736 24716 12764
rect 22741 12727 22799 12733
rect 16264 12668 18184 12696
rect 16264 12656 16270 12668
rect 19334 12656 19340 12708
rect 19392 12696 19398 12708
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 19392 12668 19533 12696
rect 19392 12656 19398 12668
rect 19521 12665 19533 12668
rect 19567 12696 19579 12699
rect 20162 12696 20168 12708
rect 19567 12668 20168 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 20162 12656 20168 12668
rect 20220 12696 20226 12708
rect 21174 12696 21180 12708
rect 20220 12668 21180 12696
rect 20220 12656 20226 12668
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 24118 12696 24124 12708
rect 24079 12668 24124 12696
rect 24118 12656 24124 12668
rect 24176 12656 24182 12708
rect 24670 12656 24676 12708
rect 24728 12696 24734 12708
rect 24771 12696 24799 12804
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 25046 12835 25104 12841
rect 25046 12801 25058 12835
rect 25092 12832 25104 12835
rect 25792 12832 25820 12872
rect 25885 12869 25897 12872
rect 25931 12869 25943 12903
rect 25885 12863 25943 12869
rect 26418 12860 26424 12912
rect 26476 12900 26482 12912
rect 27356 12909 27384 12940
rect 30009 12937 30021 12940
rect 30055 12937 30067 12971
rect 30009 12931 30067 12937
rect 27249 12903 27307 12909
rect 27249 12900 27261 12903
rect 26476 12872 27261 12900
rect 26476 12860 26482 12872
rect 27249 12869 27261 12872
rect 27295 12869 27307 12903
rect 27249 12863 27307 12869
rect 27341 12903 27399 12909
rect 27341 12869 27353 12903
rect 27387 12869 27399 12903
rect 27341 12863 27399 12869
rect 28896 12903 28954 12909
rect 28896 12869 28908 12903
rect 28942 12900 28954 12903
rect 28994 12900 29000 12912
rect 28942 12872 29000 12900
rect 28942 12869 28954 12872
rect 28896 12863 28954 12869
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 26970 12832 26976 12844
rect 25092 12804 25820 12832
rect 26931 12804 26976 12832
rect 25092 12801 25104 12804
rect 25046 12795 25104 12801
rect 25056 12764 25084 12795
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27066 12835 27124 12841
rect 27066 12801 27078 12835
rect 27112 12801 27124 12835
rect 27438 12835 27496 12841
rect 27438 12832 27450 12835
rect 27066 12795 27124 12801
rect 27356 12804 27450 12832
rect 24872 12736 25084 12764
rect 24872 12708 24900 12736
rect 25222 12724 25228 12776
rect 25280 12764 25286 12776
rect 27080 12764 27108 12795
rect 27356 12764 27384 12804
rect 27438 12801 27450 12804
rect 27484 12801 27496 12835
rect 27438 12795 27496 12801
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 28626 12832 28632 12844
rect 27672 12804 28632 12832
rect 27672 12792 27678 12804
rect 28626 12792 28632 12804
rect 28684 12792 28690 12844
rect 25280 12736 27108 12764
rect 27264 12736 27384 12764
rect 25280 12724 25286 12736
rect 27264 12708 27292 12736
rect 24728 12668 24799 12696
rect 24728 12656 24734 12668
rect 24854 12656 24860 12708
rect 24912 12656 24918 12708
rect 25038 12656 25044 12708
rect 25096 12696 25102 12708
rect 25096 12668 25912 12696
rect 25096 12656 25102 12668
rect 15286 12628 15292 12640
rect 13044 12600 14412 12628
rect 15247 12600 15292 12628
rect 13044 12588 13050 12600
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 17494 12628 17500 12640
rect 17455 12600 17500 12628
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20588 12600 21097 12628
rect 20588 12588 20594 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 21085 12591 21143 12597
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 23106 12628 23112 12640
rect 22235 12600 23112 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 24210 12588 24216 12640
rect 24268 12628 24274 12640
rect 25314 12628 25320 12640
rect 24268 12600 25320 12628
rect 24268 12588 24274 12600
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 25884 12637 25912 12668
rect 27246 12656 27252 12708
rect 27304 12656 27310 12708
rect 25869 12631 25927 12637
rect 25869 12597 25881 12631
rect 25915 12597 25927 12631
rect 25869 12591 25927 12597
rect 26053 12631 26111 12637
rect 26053 12597 26065 12631
rect 26099 12628 26111 12631
rect 26142 12628 26148 12640
rect 26099 12600 26148 12628
rect 26099 12597 26111 12600
rect 26053 12591 26111 12597
rect 26142 12588 26148 12600
rect 26200 12588 26206 12640
rect 27617 12631 27675 12637
rect 27617 12597 27629 12631
rect 27663 12628 27675 12631
rect 27890 12628 27896 12640
rect 27663 12600 27896 12628
rect 27663 12597 27675 12600
rect 27617 12591 27675 12597
rect 27890 12588 27896 12600
rect 27948 12628 27954 12640
rect 28810 12628 28816 12640
rect 27948 12600 28816 12628
rect 27948 12588 27954 12600
rect 28810 12588 28816 12600
rect 28868 12588 28874 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11388 12396 11805 12424
rect 11388 12384 11394 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 14461 12427 14519 12433
rect 12492 12396 12537 12424
rect 12492 12384 12498 12396
rect 14461 12393 14473 12427
rect 14507 12424 14519 12427
rect 14918 12424 14924 12436
rect 14507 12396 14924 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 16080 12396 17601 12424
rect 16080 12384 16086 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 17589 12387 17647 12393
rect 18800 12396 24624 12424
rect 11790 12288 11796 12300
rect 10244 12260 11796 12288
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9950 12220 9956 12232
rect 9171 12192 9956 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10244 12229 10272 12260
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 13780 12260 14105 12288
rect 13780 12248 13786 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 16206 12288 16212 12300
rect 16167 12260 16212 12288
rect 14093 12251 14151 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 10873 12183 10931 12189
rect 10888 12152 10916 12183
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13998 12220 14004 12232
rect 13587 12192 14004 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 12434 12152 12440 12164
rect 10888 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 8938 12084 8944 12096
rect 8899 12056 8944 12084
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10652 12056 10701 12084
rect 10652 12044 10658 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13044 12056 13369 12084
rect 13044 12044 13050 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 14292 12084 14320 12183
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 14884 12192 14933 12220
rect 14884 12180 14890 12192
rect 14921 12189 14933 12192
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15562 12220 15568 12232
rect 15335 12192 15568 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 16476 12223 16534 12229
rect 16476 12189 16488 12223
rect 16522 12220 16534 12223
rect 17494 12220 17500 12232
rect 16522 12192 17500 12220
rect 16522 12189 16534 12192
rect 16476 12183 16534 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18230 12220 18236 12232
rect 18191 12192 18236 12220
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 15010 12112 15016 12164
rect 15068 12152 15074 12164
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 15068 12124 15117 12152
rect 15068 12112 15074 12124
rect 15105 12121 15117 12124
rect 15151 12121 15163 12155
rect 15105 12115 15163 12121
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15243 12124 16068 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14292 12056 15485 12084
rect 13357 12047 13415 12053
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 16040 12084 16068 12124
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 18800 12152 18828 12396
rect 20622 12356 20628 12368
rect 20583 12328 20628 12356
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 22557 12359 22615 12365
rect 22557 12325 22569 12359
rect 22603 12325 22615 12359
rect 22557 12319 22615 12325
rect 23477 12359 23535 12365
rect 23477 12325 23489 12359
rect 23523 12356 23535 12359
rect 24210 12356 24216 12368
rect 23523 12328 24216 12356
rect 23523 12325 23535 12328
rect 23477 12319 23535 12325
rect 22572 12288 22600 12319
rect 24210 12316 24216 12328
rect 24268 12316 24274 12368
rect 24596 12356 24624 12396
rect 25038 12384 25044 12436
rect 25096 12424 25102 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 25096 12396 25329 12424
rect 25096 12384 25102 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 27154 12356 27160 12368
rect 24596 12328 27160 12356
rect 27154 12316 27160 12328
rect 27212 12316 27218 12368
rect 27614 12288 27620 12300
rect 22572 12260 23612 12288
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 19291 12192 21189 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 21177 12189 21189 12192
rect 21223 12220 21235 12223
rect 22738 12220 22744 12232
rect 21223 12192 22744 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 23106 12180 23112 12232
rect 23164 12220 23170 12232
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 23164 12192 23213 12220
rect 23164 12180 23170 12192
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23293 12223 23351 12229
rect 23293 12189 23305 12223
rect 23339 12220 23351 12223
rect 23382 12220 23388 12232
rect 23339 12192 23388 12220
rect 23339 12189 23351 12192
rect 23293 12183 23351 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 23584 12229 23612 12260
rect 23860 12260 26280 12288
rect 27575 12260 27620 12288
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 16172 12124 18828 12152
rect 19512 12155 19570 12161
rect 16172 12112 16178 12124
rect 19512 12121 19524 12155
rect 19558 12152 19570 12155
rect 19978 12152 19984 12164
rect 19558 12124 19984 12152
rect 19558 12121 19570 12124
rect 19512 12115 19570 12121
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20254 12112 20260 12164
rect 20312 12152 20318 12164
rect 21422 12155 21480 12161
rect 21422 12152 21434 12155
rect 20312 12124 21434 12152
rect 20312 12112 20318 12124
rect 21422 12121 21434 12124
rect 21468 12121 21480 12155
rect 22756 12152 22784 12180
rect 23474 12152 23480 12164
rect 22756 12124 23480 12152
rect 21422 12115 21480 12121
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 16298 12084 16304 12096
rect 16040 12056 16304 12084
rect 15473 12047 15531 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 18046 12084 18052 12096
rect 18007 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 21232 12056 23029 12084
rect 21232 12044 21238 12056
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 23017 12047 23075 12053
rect 23198 12044 23204 12096
rect 23256 12084 23262 12096
rect 23860 12084 23888 12260
rect 24026 12180 24032 12232
rect 24084 12220 24090 12232
rect 24486 12220 24492 12232
rect 24084 12192 24492 12220
rect 24084 12180 24090 12192
rect 24486 12180 24492 12192
rect 24544 12220 24550 12232
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 24544 12192 24685 12220
rect 24544 12180 24550 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 26142 12220 26148 12232
rect 26103 12192 26148 12220
rect 24673 12183 24731 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 26252 12229 26280 12260
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 26238 12223 26296 12229
rect 26238 12189 26250 12223
rect 26284 12189 26296 12223
rect 26238 12183 26296 12189
rect 26418 12180 26424 12232
rect 26476 12220 26482 12232
rect 26651 12223 26709 12229
rect 26476 12192 26521 12220
rect 26476 12180 26482 12192
rect 26651 12189 26663 12223
rect 26697 12220 26709 12223
rect 27246 12220 27252 12232
rect 26697 12192 27252 12220
rect 26697 12189 26709 12192
rect 26651 12183 26709 12189
rect 27246 12180 27252 12192
rect 27304 12180 27310 12232
rect 28166 12180 28172 12232
rect 28224 12220 28230 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 28224 12192 29745 12220
rect 28224 12180 28230 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 25133 12155 25191 12161
rect 25133 12121 25145 12155
rect 25179 12152 25191 12155
rect 25958 12152 25964 12164
rect 25179 12124 25964 12152
rect 25179 12121 25191 12124
rect 25133 12115 25191 12121
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 26513 12155 26571 12161
rect 26513 12121 26525 12155
rect 26559 12152 26571 12155
rect 27884 12155 27942 12161
rect 26559 12124 27752 12152
rect 26559 12121 26571 12124
rect 26513 12115 26571 12121
rect 23256 12056 23888 12084
rect 24489 12087 24547 12093
rect 23256 12044 23262 12056
rect 24489 12053 24501 12087
rect 24535 12084 24547 12087
rect 24854 12084 24860 12096
rect 24535 12056 24860 12084
rect 24535 12053 24547 12056
rect 24489 12047 24547 12053
rect 24854 12044 24860 12056
rect 24912 12084 24918 12096
rect 25222 12084 25228 12096
rect 24912 12056 25228 12084
rect 24912 12044 24918 12056
rect 25222 12044 25228 12056
rect 25280 12084 25286 12096
rect 25333 12087 25391 12093
rect 25333 12084 25345 12087
rect 25280 12056 25345 12084
rect 25280 12044 25286 12056
rect 25333 12053 25345 12056
rect 25379 12053 25391 12087
rect 25333 12047 25391 12053
rect 25501 12087 25559 12093
rect 25501 12053 25513 12087
rect 25547 12084 25559 12087
rect 25590 12084 25596 12096
rect 25547 12056 25596 12084
rect 25547 12053 25559 12056
rect 25501 12047 25559 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 26694 12044 26700 12096
rect 26752 12084 26758 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 26752 12056 26801 12084
rect 26752 12044 26758 12056
rect 26789 12053 26801 12056
rect 26835 12053 26847 12087
rect 27724 12084 27752 12124
rect 27884 12121 27896 12155
rect 27930 12152 27942 12155
rect 28442 12152 28448 12164
rect 27930 12124 28448 12152
rect 27930 12121 27942 12124
rect 27884 12115 27942 12121
rect 28442 12112 28448 12124
rect 28500 12112 28506 12164
rect 28997 12087 29055 12093
rect 28997 12084 29009 12087
rect 27724 12056 29009 12084
rect 26789 12047 26847 12053
rect 28997 12053 29009 12056
rect 29043 12053 29055 12087
rect 29546 12084 29552 12096
rect 29507 12056 29552 12084
rect 28997 12047 29055 12053
rect 29546 12044 29552 12056
rect 29604 12044 29610 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11480 11852 11897 11880
rect 11480 11840 11486 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14182 11880 14188 11892
rect 14139 11852 14188 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14182 11840 14188 11852
rect 14240 11880 14246 11892
rect 15102 11880 15108 11892
rect 14240 11852 15108 11880
rect 14240 11840 14246 11852
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15252 11852 15945 11880
rect 15252 11840 15258 11852
rect 15933 11849 15945 11852
rect 15979 11880 15991 11883
rect 17586 11880 17592 11892
rect 15979 11852 17592 11880
rect 15979 11849 15991 11852
rect 15933 11843 15991 11849
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 20254 11880 20260 11892
rect 20215 11852 20260 11880
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 20772 11852 21281 11880
rect 20772 11840 20778 11852
rect 21269 11849 21281 11852
rect 21315 11849 21327 11883
rect 21269 11843 21327 11849
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 22888 11852 23489 11880
rect 22888 11840 22894 11852
rect 23477 11849 23489 11852
rect 23523 11880 23535 11883
rect 24026 11880 24032 11892
rect 23523 11852 24032 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 25406 11880 25412 11892
rect 24136 11852 25412 11880
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 9646 11815 9704 11821
rect 9646 11812 9658 11815
rect 8996 11784 9658 11812
rect 8996 11772 9002 11784
rect 9646 11781 9658 11784
rect 9692 11781 9704 11815
rect 17212 11815 17270 11821
rect 9646 11775 9704 11781
rect 12728 11784 16988 11812
rect 7736 11747 7794 11753
rect 7736 11713 7748 11747
rect 7782 11744 7794 11747
rect 8846 11744 8852 11756
rect 7782 11716 8852 11744
rect 7782 11713 7794 11716
rect 7736 11707 7794 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 11882 11744 11888 11756
rect 11747 11716 11888 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12728 11753 12756 11784
rect 12986 11753 12992 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12308 11716 12725 11744
rect 12308 11704 12314 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12980 11744 12992 11753
rect 12947 11716 12992 11744
rect 12713 11707 12771 11713
rect 12980 11707 12992 11716
rect 12986 11704 12992 11707
rect 13044 11704 13050 11756
rect 14568 11753 14596 11784
rect 16960 11756 16988 11784
rect 17212 11781 17224 11815
rect 17258 11812 17270 11815
rect 18046 11812 18052 11824
rect 17258 11784 18052 11812
rect 17258 11781 17270 11784
rect 17212 11775 17270 11781
rect 18046 11772 18052 11784
rect 18104 11772 18110 11824
rect 20901 11815 20959 11821
rect 20901 11812 20913 11815
rect 18156 11784 20913 11812
rect 14553 11747 14611 11753
rect 14553 11713 14565 11747
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 14820 11747 14878 11753
rect 14820 11713 14832 11747
rect 14866 11744 14878 11747
rect 15286 11744 15292 11756
rect 14866 11716 15292 11744
rect 14866 11713 14878 11716
rect 14820 11707 14878 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16942 11744 16948 11756
rect 16855 11716 16948 11744
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 18156 11744 18184 11784
rect 20901 11781 20913 11784
rect 20947 11781 20959 11815
rect 20901 11775 20959 11781
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 21174 11812 21180 11824
rect 21048 11784 21180 11812
rect 21048 11772 21054 11784
rect 21131 11781 21180 11784
rect 17052 11716 18184 11744
rect 18969 11747 19027 11753
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 6604 11648 7481 11676
rect 6604 11636 6610 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 9030 11676 9036 11688
rect 8536 11648 9036 11676
rect 8536 11636 8542 11648
rect 9030 11636 9036 11648
rect 9088 11676 9094 11688
rect 9398 11676 9404 11688
rect 9088 11648 9404 11676
rect 9088 11636 9094 11648
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 10652 11648 11529 11676
rect 10652 11636 10658 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 17052 11676 17080 11716
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 15712 11648 17080 11676
rect 15712 11636 15718 11648
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18984 11676 19012 11707
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19116 11716 19625 11744
rect 19116 11704 19122 11716
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 20714 11744 20720 11756
rect 20487 11716 20720 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 21131 11747 21143 11781
rect 21177 11772 21180 11781
rect 21232 11772 21238 11824
rect 23842 11812 23848 11824
rect 21284 11784 23848 11812
rect 21177 11747 21189 11772
rect 21131 11741 21189 11747
rect 18104 11648 19012 11676
rect 18104 11636 18110 11648
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 21284 11676 21312 11784
rect 23842 11772 23848 11784
rect 23900 11772 23906 11824
rect 24136 11821 24164 11852
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 25977 11883 26035 11889
rect 25977 11880 25989 11883
rect 25516 11852 25989 11880
rect 24136 11815 24205 11821
rect 24136 11784 24159 11815
rect 24147 11781 24159 11784
rect 24193 11781 24205 11815
rect 24147 11775 24205 11781
rect 24321 11815 24379 11821
rect 24321 11781 24333 11815
rect 24367 11812 24379 11815
rect 24486 11812 24492 11824
rect 24367 11784 24492 11812
rect 24367 11781 24379 11784
rect 24321 11775 24379 11781
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 25222 11821 25228 11824
rect 24949 11815 25007 11821
rect 24949 11781 24961 11815
rect 24995 11781 25007 11815
rect 25165 11815 25228 11821
rect 25165 11812 25177 11815
rect 25135 11784 25177 11812
rect 24949 11775 25007 11781
rect 25165 11781 25177 11784
rect 25211 11781 25228 11815
rect 25165 11775 25228 11781
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22060 11716 22385 11744
rect 22060 11704 22066 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 23382 11744 23388 11756
rect 23343 11716 23388 11744
rect 22373 11707 22431 11713
rect 23382 11704 23388 11716
rect 23440 11704 23446 11756
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 19300 11648 21312 11676
rect 19300 11636 19306 11648
rect 21450 11636 21456 11688
rect 21508 11676 21514 11688
rect 22097 11679 22155 11685
rect 22097 11676 22109 11679
rect 21508 11648 22109 11676
rect 21508 11636 21514 11648
rect 22097 11645 22109 11648
rect 22143 11676 22155 11679
rect 23400 11676 23428 11704
rect 22143 11648 23428 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18966 11608 18972 11620
rect 18564 11580 18972 11608
rect 18564 11568 18570 11580
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 21100 11580 21588 11608
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 6328 11512 8861 11540
rect 6328 11500 6334 11512
rect 8849 11509 8861 11512
rect 8895 11540 8907 11543
rect 9030 11540 9036 11552
rect 8895 11512 9036 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 9640 11512 10793 11540
rect 9640 11500 9646 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17586 11540 17592 11552
rect 16632 11512 17592 11540
rect 16632 11500 16638 11512
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 17920 11512 18337 11540
rect 17920 11500 17926 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 18325 11503 18383 11509
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 18785 11543 18843 11549
rect 18785 11540 18797 11543
rect 18748 11512 18797 11540
rect 18748 11500 18754 11512
rect 18785 11509 18797 11512
rect 18831 11509 18843 11543
rect 18785 11503 18843 11509
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 21100 11549 21128 11580
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19392 11512 19441 11540
rect 19392 11500 19398 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 21085 11543 21143 11549
rect 21085 11509 21097 11543
rect 21131 11509 21143 11543
rect 21560 11540 21588 11580
rect 22002 11568 22008 11620
rect 22060 11608 22066 11620
rect 23584 11608 23612 11707
rect 24854 11676 24860 11688
rect 22060 11580 23612 11608
rect 24320 11648 24860 11676
rect 22060 11568 22066 11580
rect 22186 11540 22192 11552
rect 21560 11512 22192 11540
rect 21085 11503 21143 11509
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 24320 11549 24348 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 24964 11676 24992 11775
rect 25222 11772 25228 11775
rect 25280 11812 25286 11824
rect 25516 11812 25544 11852
rect 25977 11849 25989 11852
rect 26023 11849 26035 11883
rect 25977 11843 26035 11849
rect 27985 11883 28043 11889
rect 27985 11849 27997 11883
rect 28031 11880 28043 11883
rect 28166 11880 28172 11892
rect 28031 11852 28172 11880
rect 28031 11849 28043 11852
rect 27985 11843 28043 11849
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 28902 11840 28908 11892
rect 28960 11880 28966 11892
rect 29917 11883 29975 11889
rect 29917 11880 29929 11883
rect 28960 11852 29929 11880
rect 28960 11840 28966 11852
rect 29917 11849 29929 11852
rect 29963 11849 29975 11883
rect 29917 11843 29975 11849
rect 25280 11784 25544 11812
rect 25777 11815 25835 11821
rect 25280 11772 25286 11784
rect 25777 11781 25789 11815
rect 25823 11812 25835 11815
rect 25866 11812 25872 11824
rect 25823 11784 25872 11812
rect 25823 11781 25835 11784
rect 25777 11775 25835 11781
rect 25866 11772 25872 11784
rect 25924 11772 25930 11824
rect 27617 11815 27675 11821
rect 27617 11781 27629 11815
rect 27663 11812 27675 11815
rect 27706 11812 27712 11824
rect 27663 11784 27712 11812
rect 27663 11781 27675 11784
rect 27617 11775 27675 11781
rect 27706 11772 27712 11784
rect 27764 11772 27770 11824
rect 28804 11815 28862 11821
rect 28804 11781 28816 11815
rect 28850 11812 28862 11815
rect 29546 11812 29552 11824
rect 28850 11784 29552 11812
rect 28850 11781 28862 11784
rect 28804 11775 28862 11781
rect 29546 11772 29552 11784
rect 29604 11772 29610 11824
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26016 11716 27169 11744
rect 26016 11704 26022 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27522 11704 27528 11756
rect 27580 11744 27586 11756
rect 27801 11747 27859 11753
rect 27801 11744 27813 11747
rect 27580 11716 27813 11744
rect 27580 11704 27586 11716
rect 27801 11713 27813 11716
rect 27847 11713 27859 11747
rect 27801 11707 27859 11713
rect 28537 11747 28595 11753
rect 28537 11713 28549 11747
rect 28583 11744 28595 11747
rect 28626 11744 28632 11756
rect 28583 11716 28632 11744
rect 28583 11713 28595 11716
rect 28537 11707 28595 11713
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 28258 11676 28264 11688
rect 24964 11648 28264 11676
rect 28258 11636 28264 11648
rect 28316 11636 28322 11688
rect 24578 11568 24584 11620
rect 24636 11608 24642 11620
rect 25317 11611 25375 11617
rect 25317 11608 25329 11611
rect 24636 11580 25329 11608
rect 24636 11568 24642 11580
rect 25317 11577 25329 11580
rect 25363 11577 25375 11611
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 25317 11571 25375 11577
rect 25976 11580 26985 11608
rect 24305 11543 24363 11549
rect 24305 11509 24317 11543
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 24489 11543 24547 11549
rect 24489 11509 24501 11543
rect 24535 11540 24547 11543
rect 24946 11540 24952 11552
rect 24535 11512 24952 11540
rect 24535 11509 24547 11512
rect 24489 11503 24547 11509
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 25976 11549 26004 11580
rect 26973 11577 26985 11580
rect 27019 11577 27031 11611
rect 26973 11571 27031 11577
rect 25133 11543 25191 11549
rect 25133 11540 25145 11543
rect 25096 11512 25145 11540
rect 25096 11500 25102 11512
rect 25133 11509 25145 11512
rect 25179 11540 25191 11543
rect 25961 11543 26019 11549
rect 25961 11540 25973 11543
rect 25179 11512 25973 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 25961 11509 25973 11512
rect 26007 11509 26019 11543
rect 25961 11503 26019 11509
rect 26145 11543 26203 11549
rect 26145 11509 26157 11543
rect 26191 11540 26203 11543
rect 26510 11540 26516 11552
rect 26191 11512 26516 11540
rect 26191 11509 26203 11512
rect 26145 11503 26203 11509
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8904 11308 8953 11336
rect 8904 11296 8910 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 14737 11339 14795 11345
rect 9088 11308 14688 11336
rect 9088 11296 9094 11308
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 7708 11240 7941 11268
rect 7708 11228 7714 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 7929 11231 7987 11237
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 12989 11271 13047 11277
rect 12989 11268 13001 11271
rect 12676 11240 13001 11268
rect 12676 11228 12682 11240
rect 12989 11237 13001 11240
rect 13035 11237 13047 11271
rect 14660 11268 14688 11308
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 15470 11336 15476 11348
rect 14783 11308 15476 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 16666 11336 16672 11348
rect 15672 11308 16672 11336
rect 15672 11268 15700 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16850 11336 16856 11348
rect 16807 11308 16856 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17310 11336 17316 11348
rect 17092 11308 17316 11336
rect 17092 11296 17098 11308
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 20806 11336 20812 11348
rect 17552 11308 20812 11336
rect 17552 11296 17558 11308
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 23198 11336 23204 11348
rect 20956 11308 23204 11336
rect 20956 11296 20962 11308
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 24673 11339 24731 11345
rect 24673 11336 24685 11339
rect 23532 11308 24685 11336
rect 23532 11296 23538 11308
rect 24673 11305 24685 11308
rect 24719 11305 24731 11339
rect 24673 11299 24731 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25866 11336 25872 11348
rect 24912 11308 25872 11336
rect 24912 11296 24918 11308
rect 25866 11296 25872 11308
rect 25924 11336 25930 11348
rect 28442 11336 28448 11348
rect 25924 11308 26740 11336
rect 28403 11308 28448 11336
rect 25924 11296 25930 11308
rect 14660 11240 15700 11268
rect 15749 11271 15807 11277
rect 12989 11231 13047 11237
rect 15749 11237 15761 11271
rect 15795 11237 15807 11271
rect 17862 11268 17868 11280
rect 15749 11231 15807 11237
rect 17236 11240 17868 11268
rect 15764 11200 15792 11231
rect 14568 11172 15792 11200
rect 15948 11172 16611 11200
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 6546 11132 6552 11144
rect 4948 11104 6552 11132
rect 4948 11092 4954 11104
rect 6546 11092 6552 11104
rect 6604 11132 6610 11144
rect 8386 11132 8392 11144
rect 6604 11104 8392 11132
rect 6604 11092 6610 11104
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9456 11104 9781 11132
rect 9456 11092 9462 11104
rect 9769 11101 9781 11104
rect 9815 11132 9827 11135
rect 11606 11132 11612 11144
rect 9815 11104 11612 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14568 11141 14596 11172
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13780 11104 14381 11132
rect 13780 11092 13786 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 15194 11132 15200 11144
rect 15155 11104 15200 11132
rect 14553 11095 14611 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15562 11132 15568 11144
rect 15523 11104 15568 11132
rect 15562 11092 15568 11104
rect 15620 11132 15626 11144
rect 15948 11132 15976 11172
rect 16583 11144 16611 11172
rect 15620 11104 15976 11132
rect 15620 11092 15626 11104
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 16080 11104 16221 11132
rect 16080 11092 16086 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16209 11095 16267 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16574 11092 16580 11144
rect 16632 11141 16638 11144
rect 16632 11135 16659 11141
rect 16647 11132 16659 11135
rect 16647 11104 16725 11132
rect 16647 11101 16659 11104
rect 16632 11095 16659 11101
rect 16632 11092 16638 11095
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17236 11141 17264 11240
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 20622 11268 20628 11280
rect 20583 11240 20628 11268
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 21542 11268 21548 11280
rect 21232 11240 21548 11268
rect 21232 11228 21238 11240
rect 21542 11228 21548 11240
rect 21600 11228 21606 11280
rect 26234 11228 26240 11280
rect 26292 11268 26298 11280
rect 26292 11240 26649 11268
rect 26292 11228 26298 11240
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 17926 11172 19257 11200
rect 17926 11144 17954 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 21726 11200 21732 11212
rect 19245 11163 19303 11169
rect 20916 11172 21588 11200
rect 21687 11172 21732 11200
rect 17236 11135 17299 11141
rect 16908 11126 17080 11132
rect 16908 11104 17172 11126
rect 17236 11104 17253 11135
rect 16908 11092 16914 11104
rect 17052 11098 17172 11104
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 10042 11073 10048 11076
rect 6794 11067 6852 11073
rect 6794 11064 6806 11067
rect 6696 11036 6806 11064
rect 6696 11024 6702 11036
rect 6794 11033 6806 11036
rect 6840 11033 6852 11067
rect 10036 11064 10048 11073
rect 10003 11036 10048 11064
rect 6794 11027 6852 11033
rect 10036 11027 10048 11036
rect 10042 11024 10048 11027
rect 10100 11024 10106 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11854 11067 11912 11073
rect 11854 11064 11866 11067
rect 11020 11036 11866 11064
rect 11020 11024 11026 11036
rect 11854 11033 11866 11036
rect 11900 11033 11912 11067
rect 11854 11027 11912 11033
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 15068 11036 15393 11064
rect 15068 11024 15074 11036
rect 15381 11033 15393 11036
rect 15427 11033 15439 11067
rect 15381 11027 15439 11033
rect 15473 11067 15531 11073
rect 15473 11033 15485 11067
rect 15519 11064 15531 11067
rect 16114 11064 16120 11076
rect 15519 11036 16120 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11149 10999 11207 11005
rect 11149 10996 11161 10999
rect 10744 10968 11161 10996
rect 10744 10956 10750 10968
rect 11149 10965 11161 10968
rect 11195 10965 11207 10999
rect 15396 10996 15424 11027
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 16393 11067 16451 11073
rect 16393 11033 16405 11067
rect 16439 11033 16451 11067
rect 17144 11064 17172 11098
rect 17241 11101 17253 11104
rect 17287 11101 17299 11135
rect 17494 11132 17500 11144
rect 17455 11104 17500 11132
rect 17241 11095 17299 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 17644 11104 17689 11132
rect 17644 11092 17650 11104
rect 17862 11092 17868 11144
rect 17920 11104 17954 11144
rect 18414 11132 18420 11144
rect 18375 11104 18420 11132
rect 17920 11092 17926 11104
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 20916 11132 20944 11172
rect 21560 11144 21588 11172
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 23569 11203 23627 11209
rect 22336 11172 22784 11200
rect 22336 11160 22342 11172
rect 18564 11104 20944 11132
rect 18564 11092 18570 11104
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 21048 11104 21281 11132
rect 21048 11092 21054 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 21450 11132 21456 11144
rect 21407 11104 21456 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 22756 11141 22784 11172
rect 23569 11169 23581 11203
rect 23615 11200 23627 11203
rect 24670 11200 24676 11212
rect 23615 11172 24676 11200
rect 23615 11169 23627 11172
rect 23569 11163 23627 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 25590 11200 25596 11212
rect 25429 11172 25596 11200
rect 22741 11135 22799 11141
rect 21600 11104 21693 11132
rect 21600 11092 21606 11104
rect 22741 11101 22753 11135
rect 22787 11132 22799 11135
rect 23106 11132 23112 11144
rect 22787 11104 23112 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 23477 11135 23535 11141
rect 23477 11132 23489 11135
rect 23440 11104 23489 11132
rect 23440 11092 23446 11104
rect 23477 11101 23489 11104
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 23661 11135 23719 11141
rect 23661 11101 23673 11135
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 17405 11067 17463 11073
rect 17405 11064 17417 11067
rect 17144 11036 17417 11064
rect 16393 11027 16451 11033
rect 17405 11033 17417 11036
rect 17451 11033 17463 11067
rect 19490 11067 19548 11073
rect 19490 11064 19502 11067
rect 17405 11027 17463 11033
rect 18248 11036 19502 11064
rect 15654 10996 15660 11008
rect 15396 10968 15660 10996
rect 11149 10959 11207 10965
rect 15654 10956 15660 10968
rect 15712 10996 15718 11008
rect 16408 10996 16436 11027
rect 16850 10996 16856 11008
rect 15712 10968 16856 10996
rect 15712 10956 15718 10968
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 18248 11005 18276 11036
rect 19490 11033 19502 11036
rect 19536 11033 19548 11067
rect 19490 11027 19548 11033
rect 21082 11024 21088 11076
rect 21140 11064 21146 11076
rect 21818 11064 21824 11076
rect 21140 11036 21824 11064
rect 21140 11024 21146 11036
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 22094 11024 22100 11076
rect 22152 11064 22158 11076
rect 23676 11064 23704 11095
rect 23842 11092 23848 11144
rect 23900 11132 23906 11144
rect 25429 11141 25457 11172
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 25774 11200 25780 11212
rect 25687 11172 25780 11200
rect 25700 11141 25728 11172
rect 25774 11160 25780 11172
rect 25832 11200 25838 11212
rect 26418 11200 26424 11212
rect 25832 11172 26424 11200
rect 25832 11160 25838 11172
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 25409 11135 25467 11141
rect 23900 11104 24716 11132
rect 23900 11092 23906 11104
rect 24578 11064 24584 11076
rect 22152 11036 23704 11064
rect 24539 11036 24584 11064
rect 22152 11024 22158 11036
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 24688 11064 24716 11104
rect 25409 11101 25421 11135
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25502 11135 25560 11141
rect 25502 11101 25514 11135
rect 25548 11101 25560 11135
rect 25502 11095 25560 11101
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 25516 11064 25544 11095
rect 25866 11092 25872 11144
rect 25924 11141 25930 11144
rect 25924 11132 25932 11141
rect 26510 11132 26516 11144
rect 25924 11104 25969 11132
rect 26471 11104 26516 11132
rect 25924 11095 25932 11104
rect 25924 11092 25930 11095
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 26621 11141 26649 11240
rect 26606 11135 26664 11141
rect 26606 11101 26618 11135
rect 26652 11101 26664 11135
rect 26712 11132 26740 11308
rect 28442 11296 28448 11308
rect 28500 11296 28506 11348
rect 29086 11296 29092 11348
rect 29144 11336 29150 11348
rect 30193 11339 30251 11345
rect 30193 11336 30205 11339
rect 29144 11308 30205 11336
rect 29144 11296 29150 11308
rect 30193 11305 30205 11308
rect 30239 11305 30251 11339
rect 31478 11336 31484 11348
rect 31439 11308 31484 11336
rect 30193 11299 30251 11305
rect 31478 11296 31484 11308
rect 31536 11296 31542 11348
rect 27154 11268 27160 11280
rect 27115 11240 27160 11268
rect 27154 11228 27160 11240
rect 27212 11228 27218 11280
rect 27338 11228 27344 11280
rect 27396 11268 27402 11280
rect 27396 11240 31708 11268
rect 27396 11228 27402 11240
rect 26878 11160 26884 11212
rect 26936 11200 26942 11212
rect 26936 11172 31064 11200
rect 26936 11160 26942 11172
rect 26978 11135 27036 11141
rect 26978 11132 26990 11135
rect 26712 11104 26990 11132
rect 26606 11095 26664 11101
rect 26978 11101 26990 11104
rect 27024 11101 27036 11135
rect 26978 11095 27036 11101
rect 27617 11135 27675 11141
rect 27617 11101 27629 11135
rect 27663 11132 27675 11135
rect 27706 11132 27712 11144
rect 27663 11104 27712 11132
rect 27663 11101 27675 11104
rect 27617 11095 27675 11101
rect 27706 11092 27712 11104
rect 27764 11092 27770 11144
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 27985 11135 28043 11141
rect 27856 11104 27901 11132
rect 27856 11092 27862 11104
rect 27985 11101 27997 11135
rect 28031 11132 28043 11135
rect 28629 11135 28687 11141
rect 28629 11132 28641 11135
rect 28031 11104 28641 11132
rect 28031 11101 28043 11104
rect 27985 11095 28043 11101
rect 28629 11101 28641 11104
rect 28675 11101 28687 11135
rect 28629 11095 28687 11101
rect 28718 11092 28724 11144
rect 28776 11132 28782 11144
rect 29546 11132 29552 11144
rect 28776 11104 29552 11132
rect 28776 11092 28782 11104
rect 29546 11092 29552 11104
rect 29604 11092 29610 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29656 11104 29745 11132
rect 24688 11036 25544 11064
rect 25777 11067 25835 11073
rect 25777 11033 25789 11067
rect 25823 11064 25835 11067
rect 26234 11064 26240 11076
rect 25823 11036 26240 11064
rect 25823 11033 25835 11036
rect 25777 11027 25835 11033
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 26326 11024 26332 11076
rect 26384 11024 26390 11076
rect 26418 11024 26424 11076
rect 26476 11064 26482 11076
rect 26789 11067 26847 11073
rect 26789 11064 26801 11067
rect 26476 11036 26801 11064
rect 26476 11024 26482 11036
rect 26789 11033 26801 11036
rect 26835 11033 26847 11067
rect 26789 11027 26847 11033
rect 26881 11067 26939 11073
rect 26881 11033 26893 11067
rect 26927 11064 26939 11067
rect 26927 11036 27568 11064
rect 26927 11033 26939 11036
rect 26881 11027 26939 11033
rect 17773 10999 17831 11005
rect 17773 10996 17785 10999
rect 17092 10968 17785 10996
rect 17092 10956 17098 10968
rect 17773 10965 17785 10968
rect 17819 10965 17831 10999
rect 17773 10959 17831 10965
rect 18233 10999 18291 11005
rect 18233 10965 18245 10999
rect 18279 10965 18291 10999
rect 18233 10959 18291 10965
rect 22925 10999 22983 11005
rect 22925 10965 22937 10999
rect 22971 10996 22983 10999
rect 23198 10996 23204 11008
rect 22971 10968 23204 10996
rect 22971 10965 22983 10968
rect 22925 10959 22983 10965
rect 23198 10956 23204 10968
rect 23256 10956 23262 11008
rect 26053 10999 26111 11005
rect 26053 10965 26065 10999
rect 26099 10996 26111 10999
rect 26344 10996 26372 11024
rect 26099 10968 26372 10996
rect 27540 10996 27568 11036
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 29656 11064 29684 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 29822 11092 29828 11144
rect 29880 11132 29886 11144
rect 31036 11141 31064 11172
rect 31680 11141 31708 11240
rect 30377 11135 30435 11141
rect 30377 11132 30389 11135
rect 29880 11104 30389 11132
rect 29880 11092 29886 11104
rect 30377 11101 30389 11104
rect 30423 11101 30435 11135
rect 30377 11095 30435 11101
rect 31021 11135 31079 11141
rect 31021 11101 31033 11135
rect 31067 11101 31079 11135
rect 31021 11095 31079 11101
rect 31665 11135 31723 11141
rect 31665 11101 31677 11135
rect 31711 11101 31723 11135
rect 31665 11095 31723 11101
rect 28132 11036 29684 11064
rect 28132 11024 28138 11036
rect 28902 10996 28908 11008
rect 27540 10968 28908 10996
rect 26099 10965 26111 10968
rect 26053 10959 26111 10965
rect 28902 10956 28908 10968
rect 28960 10956 28966 11008
rect 29546 10996 29552 11008
rect 29507 10968 29552 10996
rect 29546 10956 29552 10968
rect 29604 10956 29610 11008
rect 30834 10996 30840 11008
rect 30795 10968 30840 10996
rect 30834 10956 30840 10968
rect 30892 10956 30898 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 6638 10792 6644 10804
rect 6503 10764 6644 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7469 10795 7527 10801
rect 7469 10761 7481 10795
rect 7515 10792 7527 10795
rect 9122 10792 9128 10804
rect 7515 10764 9128 10792
rect 7515 10761 7527 10764
rect 7469 10755 7527 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10008 10764 10977 10792
rect 10008 10752 10014 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11848 10764 11897 10792
rect 11848 10752 11854 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 14056 10764 14105 10792
rect 14056 10752 14062 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 18230 10792 18236 10804
rect 17175 10764 18236 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 20438 10792 20444 10804
rect 19935 10764 20444 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 21836 10764 27200 10792
rect 10612 10696 11560 10724
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7006 10656 7012 10668
rect 6687 10628 7012 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 8110 10656 8116 10668
rect 8071 10628 8116 10656
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9766 10656 9772 10668
rect 9727 10628 9772 10656
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 7098 10588 7104 10600
rect 7059 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 9876 10520 9904 10619
rect 1636 10492 9904 10520
rect 1636 10480 1642 10492
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 6788 10424 8217 10452
rect 6788 10412 6794 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8444 10424 9045 10452
rect 8444 10412 8450 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 9968 10452 9996 10619
rect 10612 10600 10640 10696
rect 11532 10665 11560 10696
rect 15010 10684 15016 10736
rect 15068 10724 15074 10736
rect 15289 10727 15347 10733
rect 15289 10724 15301 10727
rect 15068 10696 15301 10724
rect 15068 10684 15074 10696
rect 15289 10693 15301 10696
rect 15335 10693 15347 10727
rect 15289 10687 15347 10693
rect 15381 10727 15439 10733
rect 15381 10693 15393 10727
rect 15427 10724 15439 10727
rect 21836 10724 21864 10764
rect 15427 10696 21864 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 21968 10696 23521 10724
rect 21968 10684 21974 10696
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 11517 10619 11575 10625
rect 10594 10588 10600 10600
rect 10555 10560 10600 10588
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 10796 10520 10824 10619
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 15102 10656 15108 10668
rect 15063 10628 15108 10656
rect 13909 10619 13967 10625
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12713 10591 12771 10597
rect 12492 10560 12537 10588
rect 12492 10548 12498 10560
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 10183 10492 10824 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 11054 10480 11060 10532
rect 11112 10520 11118 10532
rect 12728 10520 12756 10551
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13722 10588 13728 10600
rect 12952 10560 13728 10588
rect 12952 10548 12958 10560
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13924 10588 13952 10619
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15562 10656 15568 10668
rect 15519 10628 15568 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10656 17003 10659
rect 17034 10656 17040 10668
rect 16991 10628 17040 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10656 17831 10659
rect 18138 10656 18144 10668
rect 17819 10628 18144 10656
rect 17819 10625 17831 10628
rect 17773 10619 17831 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 13924 10560 15700 10588
rect 15672 10529 15700 10560
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16632 10560 16773 10588
rect 16632 10548 16638 10560
rect 16761 10557 16773 10560
rect 16807 10557 16819 10591
rect 17862 10588 17868 10600
rect 16761 10551 16819 10557
rect 16868 10560 17868 10588
rect 11112 10492 12756 10520
rect 11112 10480 11118 10492
rect 11146 10452 11152 10464
rect 9968 10424 11152 10452
rect 9033 10415 9091 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 12728 10452 12756 10492
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10489 15715 10523
rect 15657 10483 15715 10489
rect 16868 10452 16896 10560
rect 17862 10548 17868 10560
rect 17920 10588 17926 10600
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 17920 10560 18613 10588
rect 17920 10548 17926 10560
rect 18601 10557 18613 10560
rect 18647 10557 18659 10591
rect 18601 10551 18659 10557
rect 18800 10520 18828 10619
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 19300 10628 19441 10656
rect 19300 10616 19306 10628
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 20070 10656 20076 10668
rect 19751 10628 20076 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10656 20683 10659
rect 20898 10656 20904 10668
rect 20671 10628 20904 10656
rect 20671 10625 20683 10628
rect 20625 10619 20683 10625
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 21232 10628 21281 10656
rect 21232 10616 21238 10628
rect 21269 10625 21281 10628
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 19613 10591 19671 10597
rect 19613 10557 19625 10591
rect 19659 10588 19671 10591
rect 19978 10588 19984 10600
rect 19659 10560 19984 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 21284 10588 21312 10619
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21600 10628 21833 10656
rect 21600 10616 21606 10628
rect 21821 10625 21833 10628
rect 21867 10656 21879 10659
rect 22002 10656 22008 10668
rect 21867 10628 22008 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23493 10665 23521 10696
rect 23658 10684 23664 10736
rect 23716 10724 23722 10736
rect 23716 10696 25268 10724
rect 23716 10684 23722 10696
rect 22741 10659 22799 10665
rect 22741 10656 22753 10659
rect 22388 10628 22753 10656
rect 20772 10560 21312 10588
rect 20772 10548 20778 10560
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 22388 10588 22416 10628
rect 22741 10625 22753 10628
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23478 10659 23536 10665
rect 23478 10625 23490 10659
rect 23524 10625 23536 10659
rect 23750 10656 23756 10668
rect 23711 10628 23756 10656
rect 23478 10619 23536 10625
rect 21508 10560 22416 10588
rect 22557 10591 22615 10597
rect 21508 10548 21514 10560
rect 22557 10557 22569 10591
rect 22603 10588 22615 10591
rect 23198 10588 23204 10600
rect 22603 10560 23204 10588
rect 22603 10557 22615 10560
rect 22557 10551 22615 10557
rect 23198 10548 23204 10560
rect 23256 10548 23262 10600
rect 23400 10588 23428 10619
rect 23750 10616 23756 10628
rect 23808 10616 23814 10668
rect 23891 10659 23949 10665
rect 23891 10625 23903 10659
rect 23937 10656 23949 10659
rect 24854 10656 24860 10668
rect 23937 10628 24860 10656
rect 23937 10625 23949 10628
rect 23891 10619 23949 10625
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 25240 10600 25268 10696
rect 25774 10616 25780 10668
rect 25832 10656 25838 10668
rect 25869 10659 25927 10665
rect 25869 10656 25881 10659
rect 25832 10628 25881 10656
rect 25832 10616 25838 10628
rect 25869 10625 25881 10628
rect 25915 10625 25927 10659
rect 25869 10619 25927 10625
rect 27065 10659 27123 10665
rect 27065 10625 27077 10659
rect 27111 10625 27123 10659
rect 27065 10619 27123 10625
rect 24486 10588 24492 10600
rect 23400 10560 24492 10588
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 25222 10548 25228 10600
rect 25280 10588 25286 10600
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25280 10560 25605 10588
rect 25280 10548 25286 10560
rect 25593 10557 25605 10560
rect 25639 10588 25651 10591
rect 27080 10588 27108 10619
rect 25639 10560 27108 10588
rect 27172 10588 27200 10764
rect 28902 10752 28908 10804
rect 28960 10792 28966 10804
rect 29089 10795 29147 10801
rect 29089 10792 29101 10795
rect 28960 10764 29101 10792
rect 28960 10752 28966 10764
rect 29089 10761 29101 10764
rect 29135 10761 29147 10795
rect 29089 10755 29147 10761
rect 30285 10727 30343 10733
rect 30285 10724 30297 10727
rect 27724 10696 30297 10724
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 27724 10665 27752 10696
rect 30285 10693 30297 10696
rect 30331 10693 30343 10727
rect 30285 10687 30343 10693
rect 27709 10659 27767 10665
rect 27709 10656 27721 10659
rect 27672 10628 27721 10656
rect 27672 10616 27678 10628
rect 27709 10625 27721 10628
rect 27755 10625 27767 10659
rect 27709 10619 27767 10625
rect 27976 10659 28034 10665
rect 27976 10625 27988 10659
rect 28022 10656 28034 10659
rect 29546 10656 29552 10668
rect 28022 10628 29552 10656
rect 28022 10625 28034 10628
rect 27976 10619 28034 10625
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 30101 10659 30159 10665
rect 30101 10625 30113 10659
rect 30147 10656 30159 10659
rect 30466 10656 30472 10668
rect 30147 10628 30472 10656
rect 30147 10625 30159 10628
rect 30101 10619 30159 10625
rect 30466 10616 30472 10628
rect 30524 10616 30530 10668
rect 30929 10659 30987 10665
rect 30929 10625 30941 10659
rect 30975 10625 30987 10659
rect 31570 10656 31576 10668
rect 31531 10628 31576 10656
rect 30929 10619 30987 10625
rect 27172 10560 27660 10588
rect 25639 10557 25651 10560
rect 25593 10551 25651 10557
rect 20162 10520 20168 10532
rect 18800 10492 20168 10520
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 20990 10480 20996 10532
rect 21048 10520 21054 10532
rect 21177 10523 21235 10529
rect 21177 10520 21189 10523
rect 21048 10492 21189 10520
rect 21048 10480 21054 10492
rect 21177 10489 21189 10492
rect 21223 10489 21235 10523
rect 21177 10483 21235 10489
rect 21913 10523 21971 10529
rect 21913 10489 21925 10523
rect 21959 10520 21971 10523
rect 22094 10520 22100 10532
rect 21959 10492 22100 10520
rect 21959 10489 21971 10492
rect 21913 10483 21971 10489
rect 22094 10480 22100 10492
rect 22152 10520 22158 10532
rect 22738 10520 22744 10532
rect 22152 10492 22744 10520
rect 22152 10480 22158 10492
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 22925 10523 22983 10529
rect 22925 10489 22937 10523
rect 22971 10520 22983 10523
rect 23658 10520 23664 10532
rect 22971 10492 23664 10520
rect 22971 10489 22983 10492
rect 22925 10483 22983 10489
rect 23658 10480 23664 10492
rect 23716 10480 23722 10532
rect 25041 10523 25099 10529
rect 25041 10489 25053 10523
rect 25087 10520 25099 10523
rect 27522 10520 27528 10532
rect 25087 10492 27528 10520
rect 25087 10489 25099 10492
rect 25041 10483 25099 10489
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 12728 10424 16896 10452
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 17460 10424 17601 10452
rect 17460 10412 17466 10424
rect 17589 10421 17601 10424
rect 17635 10421 17647 10455
rect 17589 10415 17647 10421
rect 18969 10455 19027 10461
rect 18969 10421 18981 10455
rect 19015 10452 19027 10455
rect 19334 10452 19340 10464
rect 19015 10424 19340 10452
rect 19015 10421 19027 10424
rect 18969 10415 19027 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 20441 10455 20499 10461
rect 20441 10421 20453 10455
rect 20487 10452 20499 10455
rect 21082 10452 21088 10464
rect 20487 10424 21088 10452
rect 20487 10421 20499 10424
rect 20441 10415 20499 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 24029 10455 24087 10461
rect 24029 10452 24041 10455
rect 23900 10424 24041 10452
rect 23900 10412 23906 10424
rect 24029 10421 24041 10424
rect 24075 10421 24087 10455
rect 24029 10415 24087 10421
rect 27062 10412 27068 10464
rect 27120 10452 27126 10464
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 27120 10424 27169 10452
rect 27120 10412 27126 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27632 10452 27660 10560
rect 28718 10548 28724 10600
rect 28776 10588 28782 10600
rect 30944 10588 30972 10619
rect 31570 10616 31576 10628
rect 31628 10616 31634 10668
rect 28776 10560 30972 10588
rect 28776 10548 28782 10560
rect 30745 10523 30803 10529
rect 30745 10489 30757 10523
rect 30791 10520 30803 10523
rect 31294 10520 31300 10532
rect 30791 10492 31300 10520
rect 30791 10489 30803 10492
rect 30745 10483 30803 10489
rect 31294 10480 31300 10492
rect 31352 10480 31358 10532
rect 30834 10452 30840 10464
rect 27632 10424 30840 10452
rect 27157 10415 27215 10421
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 31018 10412 31024 10464
rect 31076 10452 31082 10464
rect 31389 10455 31447 10461
rect 31389 10452 31401 10455
rect 31076 10424 31401 10452
rect 31076 10412 31082 10424
rect 31389 10421 31401 10424
rect 31435 10421 31447 10455
rect 31389 10415 31447 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6641 10251 6699 10257
rect 6641 10248 6653 10251
rect 6604 10220 6653 10248
rect 6604 10208 6610 10220
rect 6641 10217 6653 10220
rect 6687 10217 6699 10251
rect 6641 10211 6699 10217
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7064 10220 7941 10248
rect 7064 10208 7070 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 9999 10251 10057 10257
rect 9999 10248 10011 10251
rect 9824 10220 10011 10248
rect 9824 10208 9830 10220
rect 9999 10217 10011 10220
rect 10045 10248 10057 10251
rect 11238 10248 11244 10260
rect 10045 10220 11244 10248
rect 10045 10217 10057 10220
rect 9999 10211 10057 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 11698 10248 11704 10260
rect 11563 10220 11704 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 13906 10248 13912 10260
rect 12124 10220 13912 10248
rect 12124 10208 12130 10220
rect 13906 10208 13912 10220
rect 13964 10248 13970 10260
rect 15102 10248 15108 10260
rect 13964 10220 15108 10248
rect 13964 10208 13970 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 16942 10208 16948 10260
rect 17000 10248 17006 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 17000 10220 17509 10248
rect 17000 10208 17006 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 18693 10251 18751 10257
rect 18693 10248 18705 10251
rect 18472 10220 18705 10248
rect 18472 10208 18478 10220
rect 18693 10217 18705 10220
rect 18739 10217 18751 10251
rect 18693 10211 18751 10217
rect 19410 10251 19468 10257
rect 19410 10217 19422 10251
rect 19456 10248 19468 10251
rect 19456 10220 19656 10248
rect 19456 10217 19468 10220
rect 19410 10211 19468 10217
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 5316 10152 14473 10180
rect 5316 10140 5322 10152
rect 14461 10149 14473 10152
rect 14507 10149 14519 10183
rect 16853 10183 16911 10189
rect 16853 10180 16865 10183
rect 14461 10143 14519 10149
rect 14844 10152 16865 10180
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5184 10084 6009 10112
rect 5184 10053 5212 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7156 10084 7573 10112
rect 7156 10072 7162 10084
rect 7561 10081 7573 10084
rect 7607 10112 7619 10115
rect 11054 10112 11060 10124
rect 7607 10084 11060 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11238 10112 11244 10124
rect 11164 10084 11244 10112
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6638 10044 6644 10056
rect 6595 10016 6644 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 4982 9908 4988 9920
rect 4943 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5736 9908 5764 10007
rect 5828 9976 5856 10007
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8168 10016 9137 10044
rect 8168 10004 8174 10016
rect 9125 10013 9137 10016
rect 9171 10044 9183 10047
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9171 10016 9781 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 6914 9976 6920 9988
rect 5828 9948 6920 9976
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 9490 9976 9496 9988
rect 9355 9948 9496 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 9784 9976 9812 10007
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 11164 10053 11192 10084
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 14090 10112 14096 10124
rect 14051 10084 14096 10112
rect 14090 10072 14096 10084
rect 14148 10112 14154 10124
rect 14844 10112 14872 10152
rect 16853 10149 16865 10152
rect 16899 10149 16911 10183
rect 19058 10180 19064 10192
rect 16853 10143 16911 10149
rect 16960 10152 19064 10180
rect 15562 10112 15568 10124
rect 14148 10084 14872 10112
rect 15523 10084 15568 10112
rect 14148 10072 14154 10084
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 16960 10112 16988 10152
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 19518 10180 19524 10192
rect 19352 10152 19524 10180
rect 19352 10124 19380 10152
rect 19518 10140 19524 10152
rect 19576 10140 19582 10192
rect 19628 10180 19656 10220
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 19760 10220 19805 10248
rect 19760 10208 19766 10220
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 21600 10220 23704 10248
rect 21600 10208 21606 10220
rect 19978 10180 19984 10192
rect 19628 10152 19984 10180
rect 19978 10140 19984 10152
rect 20036 10140 20042 10192
rect 23676 10180 23704 10220
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 23845 10251 23903 10257
rect 23845 10248 23857 10251
rect 23808 10220 23857 10248
rect 23808 10208 23814 10220
rect 23845 10217 23857 10220
rect 23891 10217 23903 10251
rect 26234 10248 26240 10260
rect 23845 10211 23903 10217
rect 23952 10220 26096 10248
rect 26195 10220 26240 10248
rect 23952 10180 23980 10220
rect 23676 10152 23980 10180
rect 26068 10180 26096 10220
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 26476 10220 29776 10248
rect 26476 10208 26482 10220
rect 27338 10180 27344 10192
rect 26068 10152 27344 10180
rect 27338 10140 27344 10152
rect 27396 10140 27402 10192
rect 28813 10183 28871 10189
rect 28813 10149 28825 10183
rect 28859 10149 28871 10183
rect 28813 10143 28871 10149
rect 16172 10084 16988 10112
rect 16172 10072 16178 10084
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 17920 10084 18337 10112
rect 17920 10072 17926 10084
rect 18325 10081 18337 10084
rect 18371 10081 18383 10115
rect 19334 10112 19340 10124
rect 18325 10075 18383 10081
rect 18432 10084 19340 10112
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10744 10016 10977 10044
rect 10744 10004 10750 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11149 10007 11207 10013
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 12124 10016 12173 10044
rect 12124 10004 12130 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12492 10016 13216 10044
rect 12492 10004 12498 10016
rect 11054 9976 11060 9988
rect 9784 9948 11060 9976
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 11241 9979 11299 9985
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 11422 9976 11428 9988
rect 11287 9948 11428 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 12802 9976 12808 9988
rect 11664 9948 12808 9976
rect 11664 9936 11670 9948
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 13188 9976 13216 10016
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13964 10016 14289 10044
rect 13964 10004 13970 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15378 10044 15384 10056
rect 15335 10016 15384 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 18432 10044 18460 10084
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 20070 10112 20076 10124
rect 19659 10084 20076 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 26973 10115 27031 10121
rect 25884 10084 26832 10112
rect 16540 10016 18460 10044
rect 18509 10047 18567 10053
rect 16540 10004 16546 10016
rect 18509 10013 18521 10047
rect 18555 10013 18567 10047
rect 20990 10044 20996 10056
rect 18509 10007 18567 10013
rect 20364 10016 20996 10044
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 13188 9948 16681 9976
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16669 9939 16727 9945
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 16908 9948 17417 9976
rect 16908 9936 16914 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 18414 9936 18420 9988
rect 18472 9976 18478 9988
rect 18524 9976 18552 10007
rect 18472 9948 18552 9976
rect 19245 9979 19303 9985
rect 18472 9936 18478 9948
rect 19245 9945 19257 9979
rect 19291 9976 19303 9979
rect 20364 9976 20392 10016
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21174 10044 21180 10056
rect 21135 10016 21180 10044
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 23474 10044 23480 10056
rect 22511 10016 23480 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 23474 10004 23480 10016
rect 23532 10044 23538 10056
rect 24486 10044 24492 10056
rect 23532 10016 24492 10044
rect 23532 10004 23538 10016
rect 24486 10004 24492 10016
rect 24544 10044 24550 10056
rect 24857 10047 24915 10053
rect 24857 10044 24869 10047
rect 24544 10016 24869 10044
rect 24544 10004 24550 10016
rect 24857 10013 24869 10016
rect 24903 10013 24915 10047
rect 25884 10044 25912 10084
rect 24857 10007 24915 10013
rect 24964 10016 25912 10044
rect 19291 9948 20392 9976
rect 19291 9945 19303 9948
rect 19245 9939 19303 9945
rect 20438 9936 20444 9988
rect 20496 9976 20502 9988
rect 20533 9979 20591 9985
rect 20533 9976 20545 9979
rect 20496 9948 20545 9976
rect 20496 9936 20502 9948
rect 20533 9945 20545 9948
rect 20579 9945 20591 9979
rect 20714 9976 20720 9988
rect 20675 9948 20720 9976
rect 20533 9939 20591 9945
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 21082 9936 21088 9988
rect 21140 9976 21146 9988
rect 22710 9979 22768 9985
rect 22710 9976 22722 9979
rect 21140 9948 22722 9976
rect 21140 9936 21146 9948
rect 22710 9945 22722 9948
rect 22756 9945 22768 9979
rect 22710 9939 22768 9945
rect 23842 9936 23848 9988
rect 23900 9976 23906 9988
rect 24964 9976 24992 10016
rect 26234 10004 26240 10056
rect 26292 10044 26298 10056
rect 26697 10047 26755 10053
rect 26697 10044 26709 10047
rect 26292 10016 26709 10044
rect 26292 10004 26298 10016
rect 26697 10013 26709 10016
rect 26743 10013 26755 10047
rect 26804 10044 26832 10084
rect 26973 10081 26985 10115
rect 27019 10112 27031 10115
rect 27246 10112 27252 10124
rect 27019 10084 27252 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 27246 10072 27252 10084
rect 27304 10072 27310 10124
rect 28718 10112 28724 10124
rect 27356 10084 28724 10112
rect 27356 10044 27384 10084
rect 28718 10072 28724 10084
rect 28776 10072 28782 10124
rect 26804 10016 27384 10044
rect 26697 10007 26755 10013
rect 27706 10004 27712 10056
rect 27764 10044 27770 10056
rect 27985 10047 28043 10053
rect 27985 10044 27997 10047
rect 27764 10016 27997 10044
rect 27764 10004 27770 10016
rect 27985 10013 27997 10016
rect 28031 10044 28043 10047
rect 28828 10044 28856 10143
rect 28994 10044 29000 10056
rect 28031 10016 28856 10044
rect 28955 10016 29000 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 28994 10004 29000 10016
rect 29052 10004 29058 10056
rect 29546 10044 29552 10056
rect 29507 10016 29552 10044
rect 29546 10004 29552 10016
rect 29604 10004 29610 10056
rect 29748 10053 29776 10220
rect 30006 10072 30012 10124
rect 30064 10112 30070 10124
rect 30064 10084 31064 10112
rect 30064 10072 30070 10084
rect 29733 10047 29791 10053
rect 29733 10013 29745 10047
rect 29779 10013 29791 10047
rect 29733 10007 29791 10013
rect 29822 10004 29828 10056
rect 29880 10044 29886 10056
rect 31036 10053 31064 10084
rect 30377 10047 30435 10053
rect 30377 10044 30389 10047
rect 29880 10016 30389 10044
rect 29880 10004 29886 10016
rect 30377 10013 30389 10016
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 31021 10047 31079 10053
rect 31021 10013 31033 10047
rect 31067 10013 31079 10047
rect 31021 10007 31079 10013
rect 31386 10004 31392 10056
rect 31444 10044 31450 10056
rect 31665 10047 31723 10053
rect 31665 10044 31677 10047
rect 31444 10016 31677 10044
rect 31444 10004 31450 10016
rect 31665 10013 31677 10016
rect 31711 10013 31723 10047
rect 31665 10007 31723 10013
rect 23900 9948 24992 9976
rect 25124 9979 25182 9985
rect 23900 9936 23906 9948
rect 25124 9945 25136 9979
rect 25170 9976 25182 9979
rect 27890 9976 27896 9988
rect 25170 9948 27896 9976
rect 25170 9945 25182 9948
rect 25124 9939 25182 9945
rect 27890 9936 27896 9948
rect 27948 9936 27954 9988
rect 28166 9976 28172 9988
rect 28127 9948 28172 9976
rect 28166 9936 28172 9948
rect 28224 9936 28230 9988
rect 28353 9979 28411 9985
rect 28353 9945 28365 9979
rect 28399 9976 28411 9979
rect 30926 9976 30932 9988
rect 28399 9948 30932 9976
rect 28399 9945 28411 9948
rect 28353 9939 28411 9945
rect 30926 9936 30932 9948
rect 30984 9936 30990 9988
rect 5994 9908 6000 9920
rect 5736 9880 6000 9908
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9908 7067 9911
rect 9030 9908 9036 9920
rect 7055 9880 9036 9908
rect 7055 9877 7067 9880
rect 7009 9871 7067 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 11885 9911 11943 9917
rect 11885 9877 11897 9911
rect 11931 9908 11943 9911
rect 12066 9908 12072 9920
rect 11931 9880 12072 9908
rect 11931 9877 11943 9880
rect 11885 9871 11943 9877
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 18874 9908 18880 9920
rect 15160 9880 18880 9908
rect 15160 9868 15166 9880
rect 18874 9868 18880 9880
rect 18932 9868 18938 9920
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 20254 9908 20260 9920
rect 19392 9880 20260 9908
rect 19392 9868 19398 9880
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 26694 9868 26700 9920
rect 26752 9908 26758 9920
rect 29641 9911 29699 9917
rect 29641 9908 29653 9911
rect 26752 9880 29653 9908
rect 26752 9868 26758 9880
rect 29641 9877 29653 9880
rect 29687 9877 29699 9911
rect 30190 9908 30196 9920
rect 30151 9880 30196 9908
rect 29641 9871 29699 9877
rect 30190 9868 30196 9880
rect 30248 9868 30254 9920
rect 30282 9868 30288 9920
rect 30340 9908 30346 9920
rect 30837 9911 30895 9917
rect 30837 9908 30849 9911
rect 30340 9880 30849 9908
rect 30340 9868 30346 9880
rect 30837 9877 30849 9880
rect 30883 9877 30895 9911
rect 31478 9908 31484 9920
rect 31439 9880 31484 9908
rect 30837 9871 30895 9877
rect 31478 9868 31484 9880
rect 31536 9868 31542 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4264 9676 5028 9704
rect 4264 9636 4292 9676
rect 4890 9636 4896 9648
rect 3896 9608 4292 9636
rect 4356 9608 4896 9636
rect 3896 9577 3924 9608
rect 4356 9577 4384 9608
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5000 9636 5028 9676
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7800 9676 8217 9704
rect 7800 9664 7806 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 9490 9704 9496 9716
rect 8205 9667 8263 9673
rect 8588 9676 9496 9704
rect 8588 9648 8616 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10704 9676 12572 9704
rect 5902 9636 5908 9648
rect 5000 9608 5908 9636
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 7929 9639 7987 9645
rect 7929 9636 7941 9639
rect 6012 9608 7941 9636
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4608 9571 4666 9577
rect 4608 9537 4620 9571
rect 4654 9568 4666 9571
rect 4982 9568 4988 9580
rect 4654 9540 4988 9568
rect 4654 9537 4666 9540
rect 4608 9531 4666 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 6012 9568 6040 9608
rect 7929 9605 7941 9608
rect 7975 9605 7987 9639
rect 7929 9599 7987 9605
rect 8570 9596 8576 9648
rect 8628 9596 8634 9648
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 10704 9636 10732 9676
rect 9364 9608 10732 9636
rect 9364 9596 9370 9608
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 11793 9639 11851 9645
rect 10836 9608 10881 9636
rect 10980 9608 11744 9636
rect 10836 9596 10842 9608
rect 5408 9540 6040 9568
rect 5408 9528 5414 9540
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 6328 9540 6377 9568
rect 6328 9528 6334 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6546 9568 6552 9580
rect 6507 9540 6552 9568
rect 6365 9531 6423 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6696 9540 6929 9568
rect 6696 9528 6702 9540
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 6917 9531 6975 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 8067 9571 8125 9577
rect 8067 9537 8079 9571
rect 8113 9568 8125 9571
rect 8113 9540 8708 9568
rect 8113 9537 8125 9540
rect 8067 9531 8125 9537
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6564 9500 6592 9528
rect 6236 9472 6592 9500
rect 6825 9503 6883 9509
rect 6236 9460 6242 9472
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7742 9500 7748 9512
rect 6871 9472 7748 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 7852 9500 7880 9531
rect 8570 9500 8576 9512
rect 7852 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8680 9500 8708 9540
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 10980 9568 11008 9608
rect 8812 9540 8857 9568
rect 8956 9540 11008 9568
rect 8812 9528 8818 9540
rect 8956 9509 8984 9540
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11606 9568 11612 9580
rect 11112 9540 11612 9568
rect 11112 9528 11118 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11716 9568 11744 9608
rect 11793 9605 11805 9639
rect 11839 9636 11851 9639
rect 12342 9636 12348 9648
rect 11839 9608 12348 9636
rect 11839 9605 11851 9608
rect 11793 9599 11851 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 12544 9645 12572 9676
rect 12509 9639 12572 9645
rect 12509 9605 12521 9639
rect 12555 9608 12572 9639
rect 12636 9676 13492 9704
rect 12555 9605 12567 9608
rect 12509 9599 12567 9605
rect 12636 9568 12664 9676
rect 13464 9636 13492 9676
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 16574 9704 16580 9716
rect 13780 9676 16580 9704
rect 13780 9664 13786 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 16850 9704 16856 9716
rect 16724 9676 16856 9704
rect 16724 9664 16730 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 20993 9707 21051 9713
rect 18340 9676 20944 9704
rect 14274 9636 14280 9648
rect 13464 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 15194 9636 15200 9648
rect 14384 9608 15200 9636
rect 11716 9540 12664 9568
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 14384 9568 14412 9608
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 12860 9540 14412 9568
rect 12860 9528 12866 9540
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 15565 9571 15623 9577
rect 14516 9540 14561 9568
rect 15120 9540 15516 9568
rect 14516 9528 14522 9540
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8680 9472 8953 9500
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 9398 9500 9404 9512
rect 9359 9472 9404 9500
rect 8941 9463 8999 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9469 9735 9503
rect 12250 9500 12256 9512
rect 12211 9472 12256 9500
rect 9677 9463 9735 9469
rect 6454 9432 6460 9444
rect 5460 9404 6460 9432
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 5460 9364 5488 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 9692 9432 9720 9463
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13412 9472 14565 9500
rect 13412 9460 13418 9472
rect 14553 9469 14565 9472
rect 14599 9500 14611 9503
rect 15120 9500 15148 9540
rect 14599 9472 15148 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 15252 9472 15301 9500
rect 15252 9460 15258 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15488 9500 15516 9540
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 15654 9568 15660 9580
rect 15611 9540 15660 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 16592 9568 16620 9664
rect 18340 9636 18368 9676
rect 16776 9608 18368 9636
rect 18417 9639 18475 9645
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16592 9540 16681 9568
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16482 9500 16488 9512
rect 15488 9472 16488 9500
rect 15289 9463 15347 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 10962 9432 10968 9444
rect 9180 9404 9720 9432
rect 10923 9404 10968 9432
rect 9180 9392 9186 9404
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 14458 9432 14464 9444
rect 11532 9404 11836 9432
rect 3743 9336 5488 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5592 9336 5733 9364
rect 5592 9324 5598 9336
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 11532 9364 11560 9404
rect 9088 9336 11560 9364
rect 11808 9364 11836 9404
rect 13464 9404 14464 9432
rect 13464 9364 13492 9404
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 14829 9435 14887 9441
rect 14829 9401 14841 9435
rect 14875 9432 14887 9435
rect 16776 9432 16804 9608
rect 18417 9605 18429 9639
rect 18463 9636 18475 9639
rect 19518 9636 19524 9648
rect 18463 9608 19524 9636
rect 18463 9605 18475 9608
rect 18417 9599 18475 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 20916 9636 20944 9676
rect 20993 9673 21005 9707
rect 21039 9674 21051 9707
rect 21910 9704 21916 9716
rect 21192 9676 21916 9704
rect 21039 9673 21128 9674
rect 20993 9667 21128 9673
rect 21008 9648 21128 9667
rect 21192 9648 21220 9676
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 22428 9676 25085 9704
rect 22428 9664 22434 9676
rect 21008 9646 21088 9648
rect 20916 9608 20945 9636
rect 20917 9602 20945 9608
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17037 9571 17095 9577
rect 16908 9540 16953 9568
rect 16908 9528 16914 9540
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17681 9571 17739 9577
rect 17681 9568 17693 9571
rect 17083 9540 17693 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17681 9537 17693 9540
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 18012 9540 18153 9568
rect 18012 9528 18018 9540
rect 18141 9537 18153 9540
rect 18187 9568 18199 9571
rect 18230 9568 18236 9580
rect 18187 9540 18236 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9568 18567 9571
rect 18598 9568 18604 9580
rect 18555 9540 18604 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 17494 9460 17500 9512
rect 17552 9500 17558 9512
rect 18340 9500 18368 9531
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19869 9571 19927 9577
rect 19869 9568 19881 9571
rect 19392 9540 19881 9568
rect 19392 9528 19398 9540
rect 19869 9537 19881 9540
rect 19915 9537 19927 9571
rect 19869 9531 19927 9537
rect 20438 9528 20444 9580
rect 20496 9568 20502 9580
rect 20917 9574 21036 9602
rect 21082 9596 21088 9646
rect 21140 9596 21146 9648
rect 21174 9596 21180 9648
rect 21232 9596 21238 9648
rect 21821 9639 21879 9645
rect 21821 9605 21833 9639
rect 21867 9636 21879 9639
rect 22278 9636 22284 9648
rect 21867 9608 22284 9636
rect 21867 9605 21879 9608
rect 21821 9599 21879 9605
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 22741 9639 22799 9645
rect 22741 9605 22753 9639
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 22957 9639 23015 9645
rect 22957 9605 22969 9639
rect 23003 9636 23015 9639
rect 23750 9636 23756 9648
rect 23003 9608 23756 9636
rect 23003 9605 23015 9608
rect 22957 9599 23015 9605
rect 21008 9568 21036 9574
rect 21192 9568 21220 9596
rect 20496 9540 20852 9568
rect 21008 9540 21220 9568
rect 20496 9528 20502 9540
rect 17552 9472 18368 9500
rect 17552 9460 17558 9472
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19116 9472 19625 9500
rect 19116 9460 19122 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 20824 9500 20852 9540
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21784 9540 22017 9568
rect 21784 9528 21790 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22756 9568 22784 9599
rect 23750 9596 23756 9608
rect 23808 9596 23814 9648
rect 24670 9568 24676 9580
rect 22756 9540 24676 9568
rect 22005 9531 22063 9537
rect 24670 9528 24676 9540
rect 24728 9528 24734 9580
rect 24946 9568 24952 9580
rect 25004 9577 25010 9580
rect 25057 9577 25085 9676
rect 25222 9664 25228 9716
rect 25280 9664 25286 9716
rect 27890 9664 27896 9716
rect 27948 9704 27954 9716
rect 27985 9707 28043 9713
rect 27985 9704 27997 9707
rect 27948 9676 27997 9704
rect 27948 9664 27954 9676
rect 27985 9673 27997 9676
rect 28031 9673 28043 9707
rect 27985 9667 28043 9673
rect 30009 9707 30067 9713
rect 30009 9673 30021 9707
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 30392 9676 30880 9704
rect 25240 9577 25268 9664
rect 25317 9639 25375 9645
rect 25317 9605 25329 9639
rect 25363 9636 25375 9639
rect 25590 9636 25596 9648
rect 25363 9608 25596 9636
rect 25363 9605 25375 9608
rect 25317 9599 25375 9605
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 25682 9596 25688 9648
rect 25740 9636 25746 9648
rect 26326 9645 26332 9648
rect 26053 9639 26111 9645
rect 26053 9636 26065 9639
rect 25740 9608 26065 9636
rect 25740 9596 25746 9608
rect 26053 9605 26065 9608
rect 26099 9605 26111 9639
rect 26269 9639 26332 9645
rect 26269 9636 26281 9639
rect 26239 9608 26281 9636
rect 26053 9599 26111 9605
rect 26269 9605 26281 9608
rect 26315 9605 26332 9639
rect 26269 9599 26332 9605
rect 26326 9596 26332 9599
rect 26384 9636 26390 9648
rect 26602 9636 26608 9648
rect 26384 9608 26608 9636
rect 26384 9596 26390 9608
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 26878 9596 26884 9648
rect 26936 9636 26942 9648
rect 27062 9636 27068 9648
rect 26936 9608 27068 9636
rect 26936 9596 26942 9608
rect 27062 9596 27068 9608
rect 27120 9636 27126 9648
rect 27157 9639 27215 9645
rect 27157 9636 27169 9639
rect 27120 9608 27169 9636
rect 27120 9596 27126 9608
rect 27157 9605 27169 9608
rect 27203 9605 27215 9639
rect 27157 9599 27215 9605
rect 27249 9639 27307 9645
rect 27249 9605 27261 9639
rect 27295 9636 27307 9639
rect 30024 9636 30052 9667
rect 27295 9608 30052 9636
rect 27295 9605 27307 9608
rect 27249 9599 27307 9605
rect 30098 9596 30104 9648
rect 30156 9636 30162 9648
rect 30392 9636 30420 9676
rect 30742 9636 30748 9648
rect 30156 9608 30420 9636
rect 30484 9608 30748 9636
rect 30156 9596 30162 9608
rect 24914 9540 24952 9568
rect 24946 9528 24952 9540
rect 25004 9531 25014 9577
rect 25042 9571 25100 9577
rect 25042 9537 25054 9571
rect 25088 9537 25100 9571
rect 25042 9531 25100 9537
rect 25225 9571 25283 9577
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25414 9571 25472 9577
rect 25414 9564 25426 9571
rect 25460 9564 25472 9571
rect 25225 9531 25283 9537
rect 25004 9528 25010 9531
rect 25411 9512 25417 9564
rect 25469 9512 25475 9564
rect 26786 9528 26792 9580
rect 26844 9568 26850 9580
rect 26973 9571 27031 9577
rect 26973 9568 26985 9571
rect 26844 9540 26985 9568
rect 26844 9528 26850 9540
rect 26973 9537 26985 9540
rect 27019 9537 27031 9571
rect 27338 9568 27344 9580
rect 27299 9540 27344 9568
rect 26973 9531 27031 9537
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 28169 9571 28227 9577
rect 28169 9568 28181 9571
rect 27448 9540 28181 9568
rect 21082 9500 21088 9512
rect 20824 9472 21088 9500
rect 19613 9463 19671 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 23569 9503 23627 9509
rect 22336 9472 22381 9500
rect 22480 9472 22692 9500
rect 22336 9460 22342 9472
rect 14875 9404 16804 9432
rect 14875 9401 14887 9404
rect 14829 9395 14887 9401
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 22480 9432 22508 9472
rect 20956 9404 22508 9432
rect 22664 9432 22692 9472
rect 23569 9469 23581 9503
rect 23615 9500 23627 9503
rect 23658 9500 23664 9512
rect 23615 9472 23664 9500
rect 23615 9469 23627 9472
rect 23569 9463 23627 9469
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9500 23903 9503
rect 24854 9500 24860 9512
rect 23891 9472 24860 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 24854 9460 24860 9472
rect 24912 9460 24918 9512
rect 27448 9500 27476 9540
rect 28169 9537 28181 9540
rect 28215 9537 28227 9571
rect 28169 9531 28227 9537
rect 28896 9571 28954 9577
rect 28896 9537 28908 9571
rect 28942 9568 28954 9571
rect 30374 9568 30380 9580
rect 28942 9540 30380 9568
rect 28942 9537 28954 9540
rect 28896 9531 28954 9537
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 30484 9577 30512 9608
rect 30742 9596 30748 9608
rect 30800 9596 30806 9648
rect 30852 9636 30880 9676
rect 30852 9608 32996 9636
rect 30469 9571 30527 9577
rect 30469 9537 30481 9571
rect 30515 9537 30527 9571
rect 30469 9531 30527 9537
rect 30558 9528 30564 9580
rect 30616 9568 30622 9580
rect 30653 9571 30711 9577
rect 30653 9568 30665 9571
rect 30616 9540 30665 9568
rect 30616 9528 30622 9540
rect 30653 9537 30665 9540
rect 30699 9537 30711 9571
rect 30653 9531 30711 9537
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 26436 9472 27476 9500
rect 23109 9435 23167 9441
rect 23109 9432 23121 9435
rect 22664 9404 23121 9432
rect 20956 9392 20962 9404
rect 23109 9401 23121 9404
rect 23155 9401 23167 9435
rect 24872 9432 24900 9460
rect 25222 9432 25228 9444
rect 24872 9404 25228 9432
rect 23109 9395 23167 9401
rect 25222 9392 25228 9404
rect 25280 9392 25286 9444
rect 25774 9432 25780 9444
rect 25608 9404 25780 9432
rect 11808 9336 13492 9364
rect 13633 9367 13691 9373
rect 9088 9324 9094 9336
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 13722 9364 13728 9376
rect 13679 9336 13728 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 14918 9364 14924 9376
rect 14691 9336 14924 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 14918 9324 14924 9336
rect 14976 9364 14982 9376
rect 17218 9364 17224 9376
rect 14976 9336 17224 9364
rect 14976 9324 14982 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 18012 9336 18705 9364
rect 18012 9324 18018 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 18693 9327 18751 9333
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 22094 9364 22100 9376
rect 18932 9336 22100 9364
rect 18932 9324 18938 9336
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 22925 9367 22983 9373
rect 22244 9336 22289 9364
rect 22244 9324 22250 9336
rect 22925 9333 22937 9367
rect 22971 9364 22983 9367
rect 23014 9364 23020 9376
rect 22971 9336 23020 9364
rect 22971 9333 22983 9336
rect 22925 9327 22983 9333
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 25608 9373 25636 9404
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 26050 9392 26056 9444
rect 26108 9432 26114 9444
rect 26436 9441 26464 9472
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 28442 9500 28448 9512
rect 27672 9472 28448 9500
rect 27672 9460 27678 9472
rect 28442 9460 28448 9472
rect 28500 9500 28506 9512
rect 28629 9503 28687 9509
rect 28629 9500 28641 9503
rect 28500 9472 28641 9500
rect 28500 9460 28506 9472
rect 28629 9469 28641 9472
rect 28675 9469 28687 9503
rect 28629 9463 28687 9469
rect 29638 9460 29644 9512
rect 29696 9500 29702 9512
rect 31312 9500 31340 9531
rect 31938 9528 31944 9580
rect 31996 9568 32002 9580
rect 32968 9577 32996 9608
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 31996 9540 32321 9568
rect 31996 9528 32002 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32953 9571 33011 9577
rect 32953 9537 32965 9571
rect 32999 9537 33011 9571
rect 33594 9568 33600 9580
rect 33555 9540 33600 9568
rect 32953 9531 33011 9537
rect 33594 9528 33600 9540
rect 33652 9528 33658 9580
rect 29696 9472 31340 9500
rect 29696 9460 29702 9472
rect 26421 9435 26479 9441
rect 26108 9404 26280 9432
rect 26108 9392 26114 9404
rect 26252 9373 26280 9404
rect 26421 9401 26433 9435
rect 26467 9401 26479 9435
rect 28166 9432 28172 9444
rect 26421 9395 26479 9401
rect 27540 9404 28172 9432
rect 25593 9367 25651 9373
rect 25593 9333 25605 9367
rect 25639 9333 25651 9367
rect 25593 9327 25651 9333
rect 26237 9367 26295 9373
rect 26237 9333 26249 9367
rect 26283 9333 26295 9367
rect 26237 9327 26295 9333
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 27540 9373 27568 9404
rect 28166 9392 28172 9404
rect 28224 9392 28230 9444
rect 31478 9432 31484 9444
rect 29564 9404 31484 9432
rect 27525 9367 27583 9373
rect 27525 9364 27537 9367
rect 26844 9336 27537 9364
rect 26844 9324 26850 9336
rect 27525 9333 27537 9336
rect 27571 9333 27583 9367
rect 27525 9327 27583 9333
rect 27614 9324 27620 9376
rect 27672 9364 27678 9376
rect 29564 9364 29592 9404
rect 31478 9392 31484 9404
rect 31536 9392 31542 9444
rect 27672 9336 29592 9364
rect 30469 9367 30527 9373
rect 27672 9324 27678 9336
rect 30469 9333 30481 9367
rect 30515 9364 30527 9367
rect 30834 9364 30840 9376
rect 30515 9336 30840 9364
rect 30515 9333 30527 9336
rect 30469 9327 30527 9333
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 31110 9364 31116 9376
rect 31071 9336 31116 9364
rect 31110 9324 31116 9336
rect 31168 9324 31174 9376
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 32125 9367 32183 9373
rect 32125 9364 32137 9367
rect 31812 9336 32137 9364
rect 31812 9324 31818 9336
rect 32125 9333 32137 9336
rect 32171 9333 32183 9367
rect 32125 9327 32183 9333
rect 32490 9324 32496 9376
rect 32548 9364 32554 9376
rect 32769 9367 32827 9373
rect 32769 9364 32781 9367
rect 32548 9336 32781 9364
rect 32548 9324 32554 9336
rect 32769 9333 32781 9336
rect 32815 9333 32827 9367
rect 32769 9327 32827 9333
rect 33413 9367 33471 9373
rect 33413 9333 33425 9367
rect 33459 9364 33471 9367
rect 33502 9364 33508 9376
rect 33459 9336 33508 9364
rect 33459 9333 33471 9336
rect 33413 9327 33471 9333
rect 33502 9324 33508 9336
rect 33560 9324 33566 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3970 9160 3976 9172
rect 2516 9132 3976 9160
rect 2516 8965 2544 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7282 9160 7288 9172
rect 7055 9132 7288 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 13446 9160 13452 9172
rect 7800 9132 13452 9160
rect 7800 9120 7806 9132
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13906 9160 13912 9172
rect 13587 9132 13912 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 18506 9160 18512 9172
rect 14332 9132 18512 9160
rect 14332 9120 14338 9132
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 18598 9120 18604 9172
rect 18656 9160 18662 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18656 9132 18705 9160
rect 18656 9120 18662 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 19334 9160 19340 9172
rect 19295 9132 19340 9160
rect 18693 9123 18751 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 19794 9120 19800 9172
rect 19852 9160 19858 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19852 9132 19993 9160
rect 19852 9120 19858 9132
rect 19981 9129 19993 9132
rect 20027 9160 20039 9163
rect 20070 9160 20076 9172
rect 20027 9132 20076 9160
rect 20027 9129 20039 9132
rect 19981 9123 20039 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20990 9120 20996 9172
rect 21048 9160 21054 9172
rect 21358 9160 21364 9172
rect 21048 9132 21364 9160
rect 21048 9120 21054 9132
rect 21358 9120 21364 9132
rect 21416 9160 21422 9172
rect 22278 9160 22284 9172
rect 21416 9132 22284 9160
rect 21416 9120 21422 9132
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22428 9132 22508 9160
rect 22428 9120 22434 9132
rect 11974 9092 11980 9104
rect 5092 9064 11980 9092
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3936 8928 4077 8956
rect 3936 8916 3942 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4154 8888 4160 8900
rect 2746 8860 4160 8888
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2746 8820 2774 8860
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 4332 8891 4390 8897
rect 4332 8857 4344 8891
rect 4378 8888 4390 8891
rect 4706 8888 4712 8900
rect 4378 8860 4712 8888
rect 4378 8857 4390 8860
rect 4332 8851 4390 8857
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 2363 8792 2774 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 5092 8820 5120 9064
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 12802 9092 12808 9104
rect 12400 9064 12808 9092
rect 12400 9052 12406 9064
rect 12802 9052 12808 9064
rect 12860 9092 12866 9104
rect 13170 9092 13176 9104
rect 12860 9064 13176 9092
rect 12860 9052 12866 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 17681 9095 17739 9101
rect 17681 9061 17693 9095
rect 17727 9061 17739 9095
rect 21818 9092 21824 9104
rect 17681 9055 17739 9061
rect 18432 9064 21824 9092
rect 6730 9024 6736 9036
rect 6656 8996 6736 9024
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 6328 8928 6469 8956
rect 6328 8916 6334 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5224 8860 6224 8888
rect 5224 8848 5230 8860
rect 3476 8792 5120 8820
rect 5445 8823 5503 8829
rect 3476 8780 3482 8792
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 5718 8820 5724 8832
rect 5491 8792 5724 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 5718 8780 5724 8792
rect 5776 8820 5782 8832
rect 6086 8820 6092 8832
rect 5776 8792 6092 8820
rect 5776 8780 5782 8792
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6196 8820 6224 8860
rect 6546 8848 6552 8900
rect 6604 8888 6610 8900
rect 6656 8897 6684 8996
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 7668 8996 9321 9024
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7668 8965 7696 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 9456 8996 11928 9024
rect 9456 8984 9462 8996
rect 7653 8959 7711 8965
rect 6880 8928 7420 8956
rect 6880 8916 6886 8928
rect 6641 8891 6699 8897
rect 6641 8888 6653 8891
rect 6604 8860 6653 8888
rect 6604 8848 6610 8860
rect 6641 8857 6653 8860
rect 6687 8857 6699 8891
rect 6641 8851 6699 8857
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8857 6791 8891
rect 7392 8888 7420 8928
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 7800 8928 8401 8956
rect 7800 8916 7806 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 8389 8919 8447 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 9950 8956 9956 8968
rect 9171 8928 9956 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10318 8956 10324 8968
rect 10100 8928 10145 8956
rect 10279 8928 10324 8956
rect 10100 8916 10106 8928
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 11054 8916 11060 8968
rect 11112 8958 11118 8968
rect 11333 8959 11391 8965
rect 11112 8956 11275 8958
rect 11112 8952 11284 8956
rect 11333 8952 11345 8959
rect 11112 8930 11345 8952
rect 11112 8916 11118 8930
rect 11247 8928 11345 8930
rect 11256 8925 11345 8928
rect 11379 8925 11391 8959
rect 11514 8956 11520 8968
rect 11475 8928 11520 8956
rect 11256 8924 11391 8925
rect 11333 8919 11391 8924
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11790 8965 11796 8968
rect 11747 8959 11796 8965
rect 11747 8925 11759 8959
rect 11793 8925 11796 8959
rect 11747 8919 11796 8925
rect 11790 8916 11796 8919
rect 11848 8916 11854 8968
rect 11900 8956 11928 8996
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 12308 8996 14289 9024
rect 12308 8984 12314 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 17696 9024 17724 9055
rect 18322 9024 18328 9036
rect 17696 8996 18328 9024
rect 14277 8987 14335 8993
rect 12434 8956 12440 8968
rect 11900 8928 12440 8956
rect 12434 8916 12440 8928
rect 12492 8956 12498 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12492 8928 12541 8956
rect 12492 8916 12498 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12986 8956 12992 8968
rect 12947 8928 12992 8956
rect 12529 8919 12587 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 13096 8928 13277 8956
rect 7760 8888 7788 8916
rect 7392 8860 7788 8888
rect 8205 8891 8263 8897
rect 6733 8851 6791 8857
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8754 8888 8760 8900
rect 8251 8860 8760 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 6748 8820 6776 8851
rect 8754 8848 8760 8860
rect 8812 8888 8818 8900
rect 10060 8888 10088 8916
rect 11601 8891 11659 8897
rect 11601 8888 11613 8891
rect 8812 8860 10088 8888
rect 11532 8860 11613 8888
rect 8812 8848 8818 8860
rect 6196 8792 6776 8820
rect 7469 8823 7527 8829
rect 7469 8789 7481 8823
rect 7515 8820 7527 8823
rect 8018 8820 8024 8832
rect 7515 8792 8024 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11532 8820 11560 8860
rect 11601 8857 11613 8860
rect 11647 8857 11659 8891
rect 13096 8888 13124 8928
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13630 8956 13636 8968
rect 13403 8928 13636 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16942 8956 16948 8968
rect 16347 8928 16948 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17678 8956 17684 8968
rect 17092 8928 17684 8956
rect 17092 8916 17098 8928
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 18156 8965 18184 8996
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 18432 8965 18460 9064
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 22480 9092 22508 9132
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23014 9160 23020 9172
rect 22704 9132 23020 9160
rect 22704 9120 22710 9132
rect 23014 9120 23020 9132
rect 23072 9120 23078 9172
rect 25590 9120 25596 9172
rect 25648 9160 25654 9172
rect 25869 9163 25927 9169
rect 25869 9160 25881 9163
rect 25648 9132 25881 9160
rect 25648 9120 25654 9132
rect 25869 9129 25881 9132
rect 25915 9129 25927 9163
rect 25869 9123 25927 9129
rect 28169 9163 28227 9169
rect 28169 9129 28181 9163
rect 28215 9160 28227 9163
rect 29822 9160 29828 9172
rect 28215 9132 29828 9160
rect 28215 9129 28227 9132
rect 28169 9123 28227 9129
rect 29822 9120 29828 9132
rect 29880 9120 29886 9172
rect 30374 9120 30380 9172
rect 30432 9160 30438 9172
rect 30837 9163 30895 9169
rect 30837 9160 30849 9163
rect 30432 9132 30849 9160
rect 30432 9120 30438 9132
rect 30837 9129 30849 9132
rect 30883 9129 30895 9163
rect 30837 9123 30895 9129
rect 31110 9092 31116 9104
rect 22480 9064 23796 9092
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 19794 9024 19800 9036
rect 18932 8996 19800 9024
rect 18932 8984 18938 8996
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 20438 9024 20444 9036
rect 20272 8996 20444 9024
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 19242 8956 19248 8968
rect 18564 8928 19248 8956
rect 18564 8916 18570 8928
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19484 8928 19533 8956
rect 19484 8916 19490 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19978 8956 19984 8968
rect 19939 8928 19984 8956
rect 19521 8919 19579 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20272 8965 20300 8996
rect 20438 8984 20444 8996
rect 20496 9024 20502 9036
rect 20496 8996 22600 9024
rect 20496 8984 20502 8996
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 11601 8851 11659 8857
rect 12268 8860 13124 8888
rect 11882 8820 11888 8832
rect 10928 8792 11560 8820
rect 11843 8792 11888 8820
rect 10928 8780 10934 8792
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12268 8820 12296 8860
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 14544 8891 14602 8897
rect 13228 8860 13273 8888
rect 13228 8848 13234 8860
rect 14544 8857 14556 8891
rect 14590 8888 14602 8891
rect 16568 8891 16626 8897
rect 14590 8860 16528 8888
rect 14590 8857 14602 8860
rect 14544 8851 14602 8857
rect 12032 8792 12296 8820
rect 12345 8823 12403 8829
rect 12032 8780 12038 8792
rect 12345 8789 12357 8823
rect 12391 8820 12403 8823
rect 12894 8820 12900 8832
rect 12391 8792 12900 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 13722 8820 13728 8832
rect 13044 8792 13728 8820
rect 13044 8780 13050 8792
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 15654 8820 15660 8832
rect 15615 8792 15660 8820
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 16500 8820 16528 8860
rect 16568 8857 16580 8891
rect 16614 8888 16626 8891
rect 17494 8888 17500 8900
rect 16614 8860 17500 8888
rect 16614 8857 16626 8860
rect 16568 8851 16626 8857
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 18322 8888 18328 8900
rect 18283 8860 18328 8888
rect 18322 8848 18328 8860
rect 18380 8888 18386 8900
rect 19058 8888 19064 8900
rect 18380 8860 19064 8888
rect 18380 8848 18386 8860
rect 19058 8848 19064 8860
rect 19116 8848 19122 8900
rect 20180 8888 20208 8919
rect 20990 8916 20996 8968
rect 21048 8956 21054 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 21048 8928 21097 8956
rect 21048 8916 21054 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 21232 8928 21281 8956
rect 21232 8916 21238 8928
rect 21269 8925 21281 8928
rect 21315 8956 21327 8959
rect 22186 8956 22192 8968
rect 21315 8928 22192 8956
rect 21315 8925 21327 8928
rect 21269 8919 21327 8925
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22572 8965 22600 8996
rect 22281 8959 22339 8965
rect 22281 8925 22293 8959
rect 22327 8925 22339 8959
rect 22281 8919 22339 8925
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 20180 8860 20300 8888
rect 20272 8832 20300 8860
rect 20806 8848 20812 8900
rect 20864 8888 20870 8900
rect 21545 8891 21603 8897
rect 21545 8888 21557 8891
rect 20864 8860 21557 8888
rect 20864 8848 20870 8860
rect 21545 8857 21557 8860
rect 21591 8857 21603 8891
rect 21545 8851 21603 8857
rect 21637 8891 21695 8897
rect 21637 8857 21649 8891
rect 21683 8888 21695 8891
rect 21726 8888 21732 8900
rect 21683 8860 21732 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 21726 8848 21732 8860
rect 21784 8848 21790 8900
rect 21910 8848 21916 8900
rect 21968 8888 21974 8900
rect 22296 8888 22324 8919
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23658 8956 23664 8968
rect 23072 8928 23664 8956
rect 23072 8916 23078 8928
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 21968 8860 22324 8888
rect 22465 8891 22523 8897
rect 21968 8848 21974 8860
rect 22465 8857 22477 8891
rect 22511 8888 22523 8891
rect 22738 8888 22744 8900
rect 22511 8860 22744 8888
rect 22511 8857 22523 8860
rect 22465 8851 22523 8857
rect 22738 8848 22744 8860
rect 22796 8848 22802 8900
rect 23768 8888 23796 9064
rect 26712 9064 31116 9092
rect 24486 9024 24492 9036
rect 24447 8996 24492 9024
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 24756 8959 24814 8965
rect 24756 8925 24768 8959
rect 24802 8956 24814 8959
rect 26712 8956 26740 9064
rect 31110 9052 31116 9064
rect 31168 9052 31174 9104
rect 32214 9052 32220 9104
rect 32272 9092 32278 9104
rect 33413 9095 33471 9101
rect 33413 9092 33425 9095
rect 32272 9064 33425 9092
rect 32272 9052 32278 9064
rect 33413 9061 33425 9064
rect 33459 9061 33471 9095
rect 33413 9055 33471 9061
rect 27430 8984 27436 9036
rect 27488 9024 27494 9036
rect 28902 9024 28908 9036
rect 27488 8996 28908 9024
rect 27488 8984 27494 8996
rect 28902 8984 28908 8996
rect 28960 8984 28966 9036
rect 28994 8984 29000 9036
rect 29052 8984 29058 9036
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 29236 8996 31708 9024
rect 29236 8984 29242 8996
rect 24802 8928 26740 8956
rect 26789 8959 26847 8965
rect 24802 8925 24814 8928
rect 24756 8919 24814 8925
rect 26789 8925 26801 8959
rect 26835 8925 26847 8959
rect 26789 8919 26847 8925
rect 26804 8888 26832 8919
rect 26878 8916 26884 8968
rect 26936 8956 26942 8968
rect 26973 8959 27031 8965
rect 26973 8956 26985 8959
rect 26936 8928 26985 8956
rect 26936 8916 26942 8928
rect 26973 8925 26985 8928
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 27246 8956 27252 8968
rect 27203 8928 27252 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 27246 8916 27252 8928
rect 27304 8916 27310 8968
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27580 8928 27813 8956
rect 27580 8916 27586 8928
rect 27801 8925 27813 8928
rect 27847 8956 27859 8959
rect 27847 8928 28120 8956
rect 27847 8925 27859 8928
rect 27801 8919 27859 8925
rect 27062 8888 27068 8900
rect 23768 8860 26832 8888
rect 27023 8860 27068 8888
rect 27062 8848 27068 8860
rect 27120 8848 27126 8900
rect 27985 8891 28043 8897
rect 27985 8888 27997 8891
rect 27356 8860 27997 8888
rect 27356 8832 27384 8860
rect 27985 8857 27997 8860
rect 28031 8857 28043 8891
rect 28092 8888 28120 8928
rect 28350 8916 28356 8968
rect 28408 8956 28414 8968
rect 28721 8959 28779 8965
rect 28721 8956 28733 8959
rect 28408 8928 28733 8956
rect 28408 8916 28414 8928
rect 28721 8925 28733 8928
rect 28767 8925 28779 8959
rect 29012 8956 29040 8984
rect 28721 8919 28779 8925
rect 28828 8928 29040 8956
rect 28828 8888 28856 8928
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29420 8928 29561 8956
rect 29420 8916 29426 8928
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8956 29791 8959
rect 29914 8956 29920 8968
rect 29779 8928 29920 8956
rect 29779 8925 29791 8928
rect 29733 8919 29791 8925
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 30374 8956 30380 8968
rect 30335 8928 30380 8956
rect 30374 8916 30380 8928
rect 30432 8916 30438 8968
rect 30926 8916 30932 8968
rect 30984 8956 30990 8968
rect 31021 8959 31079 8965
rect 31021 8956 31033 8959
rect 30984 8928 31033 8956
rect 30984 8916 30990 8928
rect 31021 8925 31033 8928
rect 31067 8925 31079 8959
rect 31021 8919 31079 8925
rect 31110 8916 31116 8968
rect 31168 8956 31174 8968
rect 31680 8965 31708 8996
rect 31481 8959 31539 8965
rect 31481 8956 31493 8959
rect 31168 8928 31493 8956
rect 31168 8916 31174 8928
rect 31481 8925 31493 8928
rect 31527 8925 31539 8959
rect 31481 8919 31539 8925
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8925 31723 8959
rect 32306 8956 32312 8968
rect 32267 8928 32312 8956
rect 31665 8919 31723 8925
rect 32306 8916 32312 8928
rect 32364 8916 32370 8968
rect 32950 8956 32956 8968
rect 32911 8928 32956 8956
rect 32950 8916 32956 8928
rect 33008 8916 33014 8968
rect 33597 8959 33655 8965
rect 33597 8925 33609 8959
rect 33643 8956 33655 8959
rect 33870 8956 33876 8968
rect 33643 8928 33876 8956
rect 33643 8925 33655 8928
rect 33597 8919 33655 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 28092 8860 28856 8888
rect 27985 8851 28043 8857
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 31573 8891 31631 8897
rect 31573 8888 31585 8891
rect 29052 8860 31585 8888
rect 29052 8848 29058 8860
rect 31573 8857 31585 8860
rect 31619 8857 31631 8891
rect 31573 8851 31631 8857
rect 18690 8820 18696 8832
rect 16500 8792 18696 8820
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 20254 8780 20260 8832
rect 20312 8780 20318 8832
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8820 20499 8823
rect 20898 8820 20904 8832
rect 20487 8792 20904 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20898 8780 20904 8792
rect 20956 8820 20962 8832
rect 21174 8820 21180 8832
rect 20956 8792 21180 8820
rect 20956 8780 20962 8792
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 22097 8823 22155 8829
rect 22097 8820 22109 8823
rect 21876 8792 22109 8820
rect 21876 8780 21882 8792
rect 22097 8789 22109 8792
rect 22143 8789 22155 8823
rect 22097 8783 22155 8789
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 24394 8820 24400 8832
rect 23799 8792 24400 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 24394 8780 24400 8792
rect 24452 8820 24458 8832
rect 26234 8820 26240 8832
rect 24452 8792 26240 8820
rect 24452 8780 24458 8792
rect 26234 8780 26240 8792
rect 26292 8780 26298 8832
rect 27338 8820 27344 8832
rect 27299 8792 27344 8820
rect 27338 8780 27344 8792
rect 27396 8780 27402 8832
rect 28166 8780 28172 8832
rect 28224 8820 28230 8832
rect 29454 8820 29460 8832
rect 28224 8792 29460 8820
rect 28224 8780 28230 8792
rect 29454 8780 29460 8792
rect 29512 8780 29518 8832
rect 29638 8820 29644 8832
rect 29599 8792 29644 8820
rect 29638 8780 29644 8792
rect 29696 8780 29702 8832
rect 29822 8780 29828 8832
rect 29880 8820 29886 8832
rect 30193 8823 30251 8829
rect 30193 8820 30205 8823
rect 29880 8792 30205 8820
rect 29880 8780 29886 8792
rect 30193 8789 30205 8792
rect 30239 8789 30251 8823
rect 32122 8820 32128 8832
rect 32083 8792 32128 8820
rect 30193 8783 30251 8789
rect 32122 8780 32128 8792
rect 32180 8780 32186 8832
rect 32766 8820 32772 8832
rect 32727 8792 32772 8820
rect 32766 8780 32772 8792
rect 32824 8780 32830 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 3234 8616 3240 8628
rect 2746 8588 3240 8616
rect 2746 8548 2774 8588
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3418 8616 3424 8628
rect 3379 8588 3424 8616
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4062 8616 4068 8628
rect 4023 8588 4068 8616
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5445 8619 5503 8625
rect 4172 8588 5396 8616
rect 4172 8548 4200 8588
rect 5258 8548 5264 8560
rect 1780 8520 2774 8548
rect 2976 8520 4200 8548
rect 4264 8520 5264 8548
rect 1780 8489 1808 8520
rect 2976 8489 3004 8520
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 3602 8480 3608 8492
rect 3563 8452 3608 8480
rect 2961 8443 3019 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4264 8489 4292 8520
rect 5258 8508 5264 8520
rect 5316 8508 5322 8560
rect 5368 8548 5396 8588
rect 5445 8585 5457 8619
rect 5491 8616 5503 8619
rect 6638 8616 6644 8628
rect 5491 8588 6644 8616
rect 5491 8585 5503 8588
rect 5445 8579 5503 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7064 8588 9904 8616
rect 7064 8576 7070 8588
rect 6270 8548 6276 8560
rect 5368 8520 6276 8548
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 6546 8548 6552 8560
rect 6507 8520 6552 8548
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 8386 8548 8392 8560
rect 8036 8520 8392 8548
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4249 8443 4307 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5626 8480 5632 8492
rect 5399 8452 5632 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6086 8480 6092 8492
rect 5767 8452 6092 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6638 8480 6644 8492
rect 6599 8452 6644 8480
rect 6365 8443 6423 8449
rect 5534 8412 5540 8424
rect 5495 8384 5540 8412
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 6380 8412 6408 8443
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6822 8480 6828 8492
rect 6779 8452 6828 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7558 8480 7564 8492
rect 7519 8452 7564 8480
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8036 8489 8064 8520
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 9876 8548 9904 8588
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10008 8588 10425 8616
rect 10008 8576 10014 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 12618 8616 12624 8628
rect 11112 8588 12624 8616
rect 11112 8576 11118 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 18046 8616 18052 8628
rect 14875 8588 18052 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 19426 8616 19432 8628
rect 18156 8588 19288 8616
rect 19387 8588 19432 8616
rect 10045 8551 10103 8557
rect 9876 8520 9996 8548
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8277 8483 8335 8489
rect 8277 8480 8289 8483
rect 8168 8452 8289 8480
rect 8168 8440 8174 8452
rect 8277 8449 8289 8452
rect 8323 8449 8335 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 8277 8443 8335 8449
rect 9416 8452 9873 8480
rect 5592 8384 6408 8412
rect 5592 8372 5598 8384
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3786 8344 3792 8356
rect 2823 8316 3792 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 4706 8344 4712 8356
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 7374 8344 7380 8356
rect 5500 8316 5580 8344
rect 7335 8316 7380 8344
rect 5500 8304 5506 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 5350 8276 5356 8288
rect 3016 8248 5356 8276
rect 3016 8236 3022 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5552 8276 5580 8316
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 7892 8316 8064 8344
rect 7892 8304 7898 8316
rect 5629 8279 5687 8285
rect 5629 8276 5641 8279
rect 5552 8248 5641 8276
rect 5629 8245 5641 8248
rect 5675 8245 5687 8279
rect 5629 8239 5687 8245
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7926 8276 7932 8288
rect 6972 8248 7932 8276
rect 6972 8236 6978 8248
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8036 8276 8064 8316
rect 9030 8276 9036 8288
rect 8036 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9416 8285 9444 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 9968 8412 9996 8520
rect 10045 8517 10057 8551
rect 10091 8548 10103 8551
rect 11238 8548 11244 8560
rect 10091 8520 11244 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 11238 8508 11244 8520
rect 11296 8548 11302 8560
rect 11698 8548 11704 8560
rect 11296 8520 11704 8548
rect 11296 8508 11302 8520
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 12710 8508 12716 8560
rect 12768 8548 12774 8560
rect 12897 8551 12955 8557
rect 12897 8548 12909 8551
rect 12768 8520 12909 8548
rect 12768 8508 12774 8520
rect 12897 8517 12909 8520
rect 12943 8517 12955 8551
rect 13630 8548 13636 8560
rect 12897 8511 12955 8517
rect 13004 8520 13636 8548
rect 10134 8480 10140 8492
rect 10095 8452 10140 8480
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10318 8480 10324 8492
rect 10275 8452 10324 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10318 8440 10324 8452
rect 10376 8480 10382 8492
rect 11146 8480 11152 8492
rect 10376 8452 11152 8480
rect 10376 8440 10382 8452
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11664 8452 11805 8480
rect 11664 8440 11670 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 12621 8483 12679 8489
rect 11940 8452 12033 8480
rect 11940 8440 11946 8452
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 12802 8480 12808 8492
rect 12763 8452 12808 8480
rect 12621 8443 12679 8449
rect 11054 8412 11060 8424
rect 9968 8384 11060 8412
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11164 8412 11192 8440
rect 11900 8412 11928 8440
rect 11164 8384 11928 8412
rect 12636 8412 12664 8443
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13004 8489 13032 8520
rect 13630 8508 13636 8520
rect 13688 8508 13694 8560
rect 17304 8551 17362 8557
rect 17304 8517 17316 8551
rect 17350 8548 17362 8551
rect 17402 8548 17408 8560
rect 17350 8520 17408 8548
rect 17350 8517 17362 8520
rect 17304 8511 17362 8517
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 18156 8548 18184 8588
rect 17644 8520 18184 8548
rect 17644 8508 17650 8520
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 19153 8551 19211 8557
rect 19153 8548 19165 8551
rect 18564 8520 19165 8548
rect 18564 8508 18570 8520
rect 19153 8517 19165 8520
rect 19199 8517 19211 8551
rect 19260 8548 19288 8588
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 21818 8616 21824 8628
rect 20824 8588 21824 8616
rect 20254 8548 20260 8560
rect 19260 8520 20260 8548
rect 19153 8511 19211 8517
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 13817 8483 13875 8489
rect 13817 8480 13829 8483
rect 13596 8452 13829 8480
rect 13596 8440 13602 8452
rect 13817 8449 13829 8452
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 15194 8480 15200 8492
rect 14691 8452 15200 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 16206 8480 16212 8492
rect 15335 8452 16212 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 17000 8452 17049 8480
rect 17000 8440 17006 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8449 18935 8483
rect 19058 8480 19064 8492
rect 19019 8452 19064 8480
rect 18877 8443 18935 8449
rect 13633 8415 13691 8421
rect 12636 8384 12848 8412
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 12526 8344 12532 8356
rect 9548 8316 12532 8344
rect 9548 8304 9554 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 12820 8344 12848 8384
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 13998 8412 14004 8424
rect 13679 8384 14004 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 13998 8372 14004 8384
rect 14056 8412 14062 8424
rect 14274 8412 14280 8424
rect 14056 8384 14280 8412
rect 14056 8372 14062 8384
rect 14274 8372 14280 8384
rect 14332 8412 14338 8424
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 14332 8384 14473 8412
rect 14332 8372 14338 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 15378 8372 15384 8424
rect 15436 8412 15442 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15436 8384 15577 8412
rect 15436 8372 15442 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 18892 8412 18920 8443
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19886 8440 19892 8492
rect 19944 8480 19950 8492
rect 20824 8489 20852 8588
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 23106 8576 23112 8628
rect 23164 8576 23170 8628
rect 25038 8576 25044 8628
rect 25096 8616 25102 8628
rect 25096 8588 25141 8616
rect 25096 8576 25102 8588
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 29825 8619 29883 8625
rect 29825 8616 29837 8619
rect 28592 8588 29837 8616
rect 28592 8576 28598 8588
rect 29825 8585 29837 8588
rect 29871 8585 29883 8619
rect 30466 8616 30472 8628
rect 30427 8588 30472 8616
rect 29825 8579 29883 8585
rect 30466 8576 30472 8588
rect 30524 8576 30530 8628
rect 30650 8576 30656 8628
rect 30708 8616 30714 8628
rect 30708 8588 33456 8616
rect 30708 8576 30714 8588
rect 20993 8551 21051 8557
rect 20993 8517 21005 8551
rect 21039 8548 21051 8551
rect 21726 8548 21732 8560
rect 21039 8520 21732 8548
rect 21039 8517 21051 8520
rect 20993 8511 21051 8517
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 23014 8548 23020 8560
rect 21928 8520 23020 8548
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19944 8452 20085 8480
rect 19944 8440 19950 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 20898 8440 20904 8492
rect 20956 8480 20962 8492
rect 21111 8483 21169 8489
rect 21111 8480 21123 8483
rect 20956 8452 21001 8480
rect 20956 8440 20962 8452
rect 21100 8449 21123 8480
rect 21157 8480 21169 8483
rect 21928 8480 21956 8520
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 23124 8548 23152 8576
rect 24029 8551 24087 8557
rect 24029 8548 24041 8551
rect 23124 8520 24041 8548
rect 24029 8517 24041 8520
rect 24075 8517 24087 8551
rect 24670 8548 24676 8560
rect 24631 8520 24676 8548
rect 24029 8511 24087 8517
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 24889 8551 24947 8557
rect 24889 8517 24901 8551
rect 24935 8548 24947 8551
rect 25866 8548 25872 8560
rect 24935 8520 25872 8548
rect 24935 8517 24947 8520
rect 24889 8511 24947 8517
rect 25866 8508 25872 8520
rect 25924 8508 25930 8560
rect 26050 8508 26056 8560
rect 26108 8548 26114 8560
rect 26108 8520 27844 8548
rect 26108 8508 26114 8520
rect 21157 8452 21956 8480
rect 21157 8449 21169 8452
rect 21100 8443 21169 8449
rect 20622 8412 20628 8424
rect 18892 8384 20628 8412
rect 15565 8375 15623 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 12894 8344 12900 8356
rect 12820 8316 12900 8344
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 14090 8304 14096 8356
rect 14148 8344 14154 8356
rect 16666 8344 16672 8356
rect 14148 8316 16672 8344
rect 14148 8304 14154 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 17972 8316 18828 8344
rect 9401 8279 9459 8285
rect 9401 8276 9413 8279
rect 9364 8248 9413 8276
rect 9364 8236 9370 8248
rect 9401 8245 9413 8248
rect 9447 8245 9459 8279
rect 9401 8239 9459 8245
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11112 8248 12081 8276
rect 11112 8236 11118 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 13173 8279 13231 8285
rect 13173 8276 13185 8279
rect 12492 8248 13185 8276
rect 12492 8236 12498 8248
rect 13173 8245 13185 8248
rect 13219 8245 13231 8279
rect 13998 8276 14004 8288
rect 13959 8248 14004 8276
rect 13173 8239 13231 8245
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 17972 8276 18000 8316
rect 14516 8248 18000 8276
rect 14516 8236 14522 8248
rect 18230 8236 18236 8288
rect 18288 8276 18294 8288
rect 18417 8279 18475 8285
rect 18417 8276 18429 8279
rect 18288 8248 18429 8276
rect 18288 8236 18294 8248
rect 18417 8245 18429 8248
rect 18463 8245 18475 8279
rect 18800 8276 18828 8316
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 19889 8347 19947 8353
rect 19889 8344 19901 8347
rect 18932 8316 19901 8344
rect 18932 8304 18938 8316
rect 19889 8313 19901 8316
rect 19935 8313 19947 8347
rect 19889 8307 19947 8313
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 21100 8344 21128 8443
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 23109 8483 23167 8489
rect 22060 8452 22105 8480
rect 22060 8440 22066 8452
rect 23109 8449 23121 8483
rect 23155 8480 23167 8483
rect 23474 8480 23480 8492
rect 23155 8452 23480 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 23474 8440 23480 8452
rect 23532 8440 23538 8492
rect 24118 8440 24124 8492
rect 24176 8480 24182 8492
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 24176 8452 25697 8480
rect 24176 8440 24182 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 26234 8480 26240 8492
rect 26195 8452 26240 8480
rect 25685 8443 25743 8449
rect 26234 8440 26240 8452
rect 26292 8440 26298 8492
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8449 27031 8483
rect 27154 8480 27160 8492
rect 27115 8452 27160 8480
rect 26973 8443 27031 8449
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21315 8384 21404 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 20036 8316 21128 8344
rect 20036 8304 20042 8316
rect 21376 8288 21404 8384
rect 23014 8372 23020 8424
rect 23072 8412 23078 8424
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 23072 8384 23213 8412
rect 23072 8372 23078 8384
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 26988 8412 27016 8443
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27816 8489 27844 8520
rect 27890 8508 27896 8560
rect 27948 8548 27954 8560
rect 27948 8520 28028 8548
rect 27948 8508 27954 8520
rect 28000 8489 28028 8520
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 30377 8551 30435 8557
rect 30377 8548 30389 8551
rect 28960 8520 30389 8548
rect 28960 8508 28966 8520
rect 30377 8517 30389 8520
rect 30423 8517 30435 8551
rect 30377 8511 30435 8517
rect 30484 8520 31754 8548
rect 27801 8483 27859 8489
rect 27801 8449 27813 8483
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 27985 8483 28043 8489
rect 27985 8449 27997 8483
rect 28031 8449 28043 8483
rect 28442 8480 28448 8492
rect 28403 8452 28448 8480
rect 27985 8443 28043 8449
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 28712 8483 28770 8489
rect 28712 8449 28724 8483
rect 28758 8480 28770 8483
rect 30190 8480 30196 8492
rect 28758 8452 30196 8480
rect 28758 8449 28770 8452
rect 28712 8443 28770 8449
rect 30190 8440 30196 8452
rect 30248 8440 30254 8492
rect 27062 8412 27068 8424
rect 23339 8384 23428 8412
rect 26975 8384 27068 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 22646 8304 22652 8356
rect 22704 8344 22710 8356
rect 23400 8344 23428 8384
rect 27062 8372 27068 8384
rect 27120 8412 27126 8424
rect 27522 8412 27528 8424
rect 27120 8384 27528 8412
rect 27120 8372 27126 8384
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 27893 8415 27951 8421
rect 27893 8412 27905 8415
rect 27580 8384 27905 8412
rect 27580 8372 27586 8384
rect 27893 8381 27905 8384
rect 27939 8381 27951 8415
rect 29822 8412 29828 8424
rect 27893 8375 27951 8381
rect 29472 8384 29828 8412
rect 24210 8344 24216 8356
rect 22704 8316 23336 8344
rect 23400 8316 24216 8344
rect 22704 8304 22710 8316
rect 20438 8276 20444 8288
rect 18800 8248 20444 8276
rect 18417 8239 18475 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 20625 8279 20683 8285
rect 20625 8245 20637 8279
rect 20671 8276 20683 8279
rect 20714 8276 20720 8288
rect 20671 8248 20720 8276
rect 20671 8245 20683 8248
rect 20625 8239 20683 8245
rect 20714 8236 20720 8248
rect 20772 8276 20778 8288
rect 21266 8276 21272 8288
rect 20772 8248 21272 8276
rect 20772 8236 20778 8248
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 21358 8236 21364 8288
rect 21416 8236 21422 8288
rect 21818 8276 21824 8288
rect 21779 8248 21824 8276
rect 21818 8236 21824 8248
rect 21876 8236 21882 8288
rect 22741 8279 22799 8285
rect 22741 8245 22753 8279
rect 22787 8276 22799 8279
rect 23014 8276 23020 8288
rect 22787 8248 23020 8276
rect 22787 8245 22799 8248
rect 22741 8239 22799 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 23308 8276 23336 8316
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 24946 8304 24952 8356
rect 25004 8344 25010 8356
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 25004 8316 25513 8344
rect 25004 8304 25010 8316
rect 25501 8313 25513 8316
rect 25547 8313 25559 8347
rect 25501 8307 25559 8313
rect 27341 8347 27399 8353
rect 27341 8313 27353 8347
rect 27387 8344 27399 8347
rect 28074 8344 28080 8356
rect 27387 8316 28080 8344
rect 27387 8313 27399 8316
rect 27341 8307 27399 8313
rect 28074 8304 28080 8316
rect 28132 8304 28138 8356
rect 29472 8344 29500 8384
rect 29822 8372 29828 8384
rect 29880 8372 29886 8424
rect 29380 8316 29500 8344
rect 24857 8279 24915 8285
rect 24857 8276 24869 8279
rect 23308 8248 24869 8276
rect 24857 8245 24869 8248
rect 24903 8276 24915 8279
rect 26050 8276 26056 8288
rect 24903 8248 26056 8276
rect 24903 8245 24915 8248
rect 24857 8239 24915 8245
rect 26050 8236 26056 8248
rect 26108 8236 26114 8288
rect 26329 8279 26387 8285
rect 26329 8245 26341 8279
rect 26375 8276 26387 8279
rect 28166 8276 28172 8288
rect 26375 8248 28172 8276
rect 26375 8245 26387 8248
rect 26329 8239 26387 8245
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 28810 8236 28816 8288
rect 28868 8276 28874 8288
rect 29380 8276 29408 8316
rect 29730 8304 29736 8356
rect 29788 8344 29794 8356
rect 30484 8344 30512 8520
rect 30650 8440 30656 8492
rect 30708 8480 30714 8492
rect 31205 8483 31263 8489
rect 31205 8480 31217 8483
rect 30708 8452 31217 8480
rect 30708 8440 30714 8452
rect 31205 8449 31217 8452
rect 31251 8449 31263 8483
rect 31726 8480 31754 8520
rect 33428 8492 33456 8588
rect 33778 8576 33784 8628
rect 33836 8616 33842 8628
rect 34425 8619 34483 8625
rect 34425 8616 34437 8619
rect 33836 8588 34437 8616
rect 33836 8576 33842 8588
rect 34425 8585 34437 8588
rect 34471 8585 34483 8619
rect 34425 8579 34483 8585
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31726 8452 32321 8480
rect 31205 8443 31263 8449
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 33226 8440 33232 8492
rect 33284 8480 33290 8492
rect 33321 8483 33379 8489
rect 33321 8480 33333 8483
rect 33284 8452 33333 8480
rect 33284 8440 33290 8452
rect 33321 8449 33333 8452
rect 33367 8449 33379 8483
rect 33321 8443 33379 8449
rect 33410 8440 33416 8492
rect 33468 8480 33474 8492
rect 33965 8483 34023 8489
rect 33965 8480 33977 8483
rect 33468 8452 33977 8480
rect 33468 8440 33474 8452
rect 33965 8449 33977 8452
rect 34011 8480 34023 8483
rect 34609 8483 34667 8489
rect 34609 8480 34621 8483
rect 34011 8452 34621 8480
rect 34011 8449 34023 8452
rect 33965 8443 34023 8449
rect 34609 8449 34621 8452
rect 34655 8449 34667 8483
rect 34609 8443 34667 8449
rect 35253 8483 35311 8489
rect 35253 8449 35265 8483
rect 35299 8480 35311 8483
rect 35342 8480 35348 8492
rect 35299 8452 35348 8480
rect 35299 8449 35311 8452
rect 35253 8443 35311 8449
rect 35342 8440 35348 8452
rect 35400 8440 35406 8492
rect 29788 8316 30512 8344
rect 30576 8384 32168 8412
rect 29788 8304 29794 8316
rect 28868 8248 29408 8276
rect 28868 8236 28874 8248
rect 30190 8236 30196 8288
rect 30248 8276 30254 8288
rect 30576 8276 30604 8384
rect 31021 8347 31079 8353
rect 31021 8313 31033 8347
rect 31067 8344 31079 8347
rect 31846 8344 31852 8356
rect 31067 8316 31852 8344
rect 31067 8313 31079 8316
rect 31021 8307 31079 8313
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 32140 8353 32168 8384
rect 32125 8347 32183 8353
rect 32125 8313 32137 8347
rect 32171 8313 32183 8347
rect 32125 8307 32183 8313
rect 33781 8347 33839 8353
rect 33781 8313 33793 8347
rect 33827 8344 33839 8347
rect 34054 8344 34060 8356
rect 33827 8316 34060 8344
rect 33827 8313 33839 8316
rect 33781 8307 33839 8313
rect 34054 8304 34060 8316
rect 34112 8304 34118 8356
rect 34514 8304 34520 8356
rect 34572 8344 34578 8356
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34572 8316 35081 8344
rect 34572 8304 34578 8316
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 30248 8248 30604 8276
rect 30248 8236 30254 8248
rect 32858 8236 32864 8288
rect 32916 8276 32922 8288
rect 33137 8279 33195 8285
rect 33137 8276 33149 8279
rect 32916 8248 33149 8276
rect 32916 8236 32922 8248
rect 33137 8245 33149 8248
rect 33183 8245 33195 8279
rect 33137 8239 33195 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 4948 8044 5457 8072
rect 4948 8032 4954 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6362 8072 6368 8084
rect 6052 8044 6368 8072
rect 6052 8032 6058 8044
rect 6362 8032 6368 8044
rect 6420 8072 6426 8084
rect 7834 8072 7840 8084
rect 6420 8044 7840 8072
rect 6420 8032 6426 8044
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 9766 8072 9772 8084
rect 7984 8044 9772 8072
rect 7984 8032 7990 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 11146 8072 11152 8084
rect 9876 8044 11152 8072
rect 9876 8004 9904 8044
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 11256 8044 14105 8072
rect 4632 7976 9904 8004
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1360 7840 1961 7868
rect 1360 7828 1366 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2866 7868 2872 7880
rect 2639 7840 2872 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3510 7868 3516 7880
rect 3283 7840 3516 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4522 7868 4528 7880
rect 4019 7840 4528 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4632 7877 4660 7976
rect 5074 7936 5080 7948
rect 5035 7908 5080 7936
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5994 7936 6000 7948
rect 5184 7908 6000 7936
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 5184 7800 5212 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7300 7908 8125 7936
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 2424 7772 5212 7800
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 1946 7732 1952 7744
rect 1811 7704 1952 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2424 7741 2452 7772
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7701 2467 7735
rect 2409 7695 2467 7701
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3384 7704 3801 7732
rect 3384 7692 3390 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 5074 7732 5080 7744
rect 4479 7704 5080 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5276 7732 5304 7831
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 5776 7840 5917 7868
rect 5776 7828 5782 7840
rect 5905 7837 5917 7840
rect 5951 7837 5963 7871
rect 6181 7871 6239 7877
rect 6181 7868 6193 7871
rect 5905 7831 5963 7837
rect 6012 7840 6193 7868
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 6012 7800 6040 7840
rect 6181 7837 6193 7840
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 6822 7868 6828 7880
rect 6319 7840 6828 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7300 7877 7328 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7834 7868 7840 7880
rect 7795 7840 7840 7868
rect 7285 7831 7343 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 5408 7772 6040 7800
rect 6089 7803 6147 7809
rect 5408 7760 5414 7772
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 6546 7800 6552 7812
rect 6135 7772 6552 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 6546 7760 6552 7772
rect 6604 7800 6610 7812
rect 7944 7800 7972 7831
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 8996 7840 9873 7868
rect 8996 7828 9002 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 8386 7800 8392 7812
rect 6604 7772 7328 7800
rect 7944 7772 8392 7800
rect 6604 7760 6610 7772
rect 7300 7744 7328 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 9217 7803 9275 7809
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 10128 7803 10186 7809
rect 9263 7772 9674 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5276 7704 6469 7732
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 6457 7695 6515 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 6972 7704 7113 7732
rect 6972 7692 6978 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9180 7704 9321 7732
rect 9180 7692 9186 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9646 7732 9674 7772
rect 10128 7769 10140 7803
rect 10174 7800 10186 7803
rect 11256 7800 11284 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16853 8075 16911 8081
rect 16853 8072 16865 8075
rect 16264 8044 16865 8072
rect 16264 8032 16270 8044
rect 16853 8041 16865 8044
rect 16899 8041 16911 8075
rect 18138 8072 18144 8084
rect 18099 8044 18144 8072
rect 16853 8035 16911 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 20162 8072 20168 8084
rect 19843 8044 20168 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 21358 8032 21364 8084
rect 21416 8072 21422 8084
rect 21453 8075 21511 8081
rect 21453 8072 21465 8075
rect 21416 8044 21465 8072
rect 21416 8032 21422 8044
rect 21453 8041 21465 8044
rect 21499 8041 21511 8075
rect 23474 8072 23480 8084
rect 21453 8035 21511 8041
rect 22066 8044 23051 8072
rect 23435 8044 23480 8072
rect 15378 8004 15384 8016
rect 12728 7976 14596 8004
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 12526 7868 12532 7880
rect 11747 7840 12532 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 10174 7772 11284 7800
rect 11968 7803 12026 7809
rect 10174 7769 10186 7772
rect 10128 7763 10186 7769
rect 11968 7769 11980 7803
rect 12014 7800 12026 7803
rect 12728 7800 12756 7976
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 14476 7800 14504 7828
rect 12014 7772 12756 7800
rect 12820 7772 14504 7800
rect 14568 7800 14596 7976
rect 14752 7976 15384 8004
rect 14752 7945 14780 7976
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 16022 7964 16028 8016
rect 16080 8004 16086 8016
rect 22066 8004 22094 8044
rect 16080 7976 22094 8004
rect 23023 8004 23051 8044
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 26237 8075 26295 8081
rect 26237 8072 26249 8075
rect 24636 8044 26249 8072
rect 24636 8032 24642 8044
rect 26237 8041 26249 8044
rect 26283 8041 26295 8075
rect 26237 8035 26295 8041
rect 27246 8032 27252 8084
rect 27304 8072 27310 8084
rect 27522 8072 27528 8084
rect 27304 8044 27528 8072
rect 27304 8032 27310 8044
rect 27522 8032 27528 8044
rect 27580 8072 27586 8084
rect 29178 8072 29184 8084
rect 27580 8044 29184 8072
rect 27580 8032 27586 8044
rect 29178 8032 29184 8044
rect 29236 8032 29242 8084
rect 31110 8072 31116 8084
rect 30392 8044 31116 8072
rect 24118 8004 24124 8016
rect 23023 7976 24124 8004
rect 16080 7964 16086 7976
rect 24118 7964 24124 7976
rect 24176 7964 24182 8016
rect 25041 8007 25099 8013
rect 25041 7973 25053 8007
rect 25087 8004 25099 8007
rect 25130 8004 25136 8016
rect 25087 7976 25136 8004
rect 25087 7973 25099 7976
rect 25041 7967 25099 7973
rect 25130 7964 25136 7976
rect 25188 7964 25194 8016
rect 28626 7964 28632 8016
rect 28684 8004 28690 8016
rect 30392 8004 30420 8044
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 33042 8032 33048 8084
rect 33100 8072 33106 8084
rect 33781 8075 33839 8081
rect 33781 8072 33793 8075
rect 33100 8044 33793 8072
rect 33100 8032 33106 8044
rect 33781 8041 33793 8044
rect 33827 8041 33839 8075
rect 33781 8035 33839 8041
rect 32122 8004 32128 8016
rect 28684 7976 30420 8004
rect 31772 7976 32128 8004
rect 28684 7964 28690 7976
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 15344 7908 16313 7936
rect 15344 7896 15350 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 21818 7936 21824 7948
rect 16301 7899 16359 7905
rect 16776 7908 21824 7936
rect 15010 7868 15016 7880
rect 14971 7840 15016 7868
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15988 7840 16037 7868
rect 15988 7828 15994 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16206 7868 16212 7880
rect 16167 7840 16212 7868
rect 16025 7831 16083 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16776 7800 16804 7908
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 23934 7936 23940 7948
rect 23716 7908 23940 7936
rect 23716 7896 23722 7908
rect 23934 7896 23940 7908
rect 23992 7896 23998 7948
rect 27065 7939 27123 7945
rect 27065 7936 27077 7939
rect 24136 7908 27077 7936
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17586 7868 17592 7880
rect 17175 7840 17592 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17954 7868 17960 7880
rect 17915 7840 17960 7868
rect 17773 7831 17831 7837
rect 14568 7772 16804 7800
rect 12014 7769 12026 7772
rect 11968 7763 12026 7769
rect 10962 7732 10968 7744
rect 9646 7704 10968 7732
rect 9309 7695 9367 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11238 7732 11244 7744
rect 11199 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7732 11302 7744
rect 11514 7732 11520 7744
rect 11296 7704 11520 7732
rect 11296 7692 11302 7704
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12820 7732 12848 7772
rect 16850 7760 16856 7812
rect 16908 7800 16914 7812
rect 17788 7800 17816 7831
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18984 7840 19257 7868
rect 17862 7800 17868 7812
rect 16908 7772 16953 7800
rect 17788 7772 17868 7800
rect 16908 7760 16914 7772
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 11940 7704 12848 7732
rect 11940 7692 11946 7704
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 13081 7735 13139 7741
rect 13081 7732 13093 7735
rect 12952 7704 13093 7732
rect 12952 7692 12958 7704
rect 13081 7701 13093 7704
rect 13127 7701 13139 7735
rect 13081 7695 13139 7701
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 15562 7732 15568 7744
rect 14516 7704 15568 7732
rect 14516 7692 14522 7704
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 17034 7732 17040 7744
rect 16995 7704 17040 7732
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 18984 7732 19012 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19392 7840 19625 7868
rect 19392 7828 19398 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20070 7868 20076 7880
rect 19944 7840 20076 7868
rect 19944 7828 19950 7840
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20680 7840 20913 7868
rect 20680 7828 20686 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21324 7840 21373 7868
rect 21324 7828 21330 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 22094 7868 22100 7880
rect 22055 7840 22100 7868
rect 21361 7831 21419 7837
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 24136 7868 24164 7908
rect 27065 7905 27077 7908
rect 27111 7936 27123 7939
rect 27111 7908 27660 7936
rect 27111 7905 27123 7908
rect 27065 7899 27123 7905
rect 22296 7840 24164 7868
rect 19058 7760 19064 7812
rect 19116 7800 19122 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 19116 7772 19441 7800
rect 19116 7760 19122 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 19429 7763 19487 7769
rect 19521 7803 19579 7809
rect 19521 7769 19533 7803
rect 19567 7800 19579 7803
rect 20254 7800 20260 7812
rect 19567 7772 20260 7800
rect 19567 7769 19579 7772
rect 19521 7763 19579 7769
rect 20254 7760 20260 7772
rect 20312 7760 20318 7812
rect 20806 7800 20812 7812
rect 20640 7772 20812 7800
rect 20640 7732 20668 7772
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 21634 7760 21640 7812
rect 21692 7800 21698 7812
rect 22002 7800 22008 7812
rect 21692 7772 22008 7800
rect 21692 7760 21698 7772
rect 22002 7760 22008 7772
rect 22060 7800 22066 7812
rect 22296 7800 22324 7840
rect 24210 7828 24216 7880
rect 24268 7868 24274 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24268 7840 24869 7868
rect 24268 7828 24274 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 26145 7871 26203 7877
rect 26145 7837 26157 7871
rect 26191 7868 26203 7871
rect 27430 7868 27436 7880
rect 26191 7840 27436 7868
rect 26191 7837 26203 7840
rect 26145 7831 26203 7837
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 27525 7871 27583 7877
rect 27525 7837 27537 7871
rect 27571 7837 27583 7871
rect 27632 7868 27660 7908
rect 28534 7896 28540 7948
rect 28592 7936 28598 7948
rect 29178 7936 29184 7948
rect 28592 7908 29184 7936
rect 28592 7896 28598 7908
rect 29178 7896 29184 7908
rect 29236 7936 29242 7948
rect 30469 7939 30527 7945
rect 30469 7936 30481 7939
rect 29236 7908 30481 7936
rect 29236 7896 29242 7908
rect 30469 7905 30481 7908
rect 30515 7905 30527 7939
rect 30469 7899 30527 7905
rect 27792 7871 27850 7877
rect 27632 7840 27752 7868
rect 27525 7831 27583 7837
rect 22060 7772 22324 7800
rect 22364 7803 22422 7809
rect 22060 7760 22066 7772
rect 22364 7769 22376 7803
rect 22410 7800 22422 7803
rect 24670 7800 24676 7812
rect 22410 7772 24676 7800
rect 22410 7769 22422 7772
rect 22364 7763 22422 7769
rect 24670 7760 24676 7772
rect 24728 7760 24734 7812
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 26418 7800 26424 7812
rect 26292 7772 26424 7800
rect 26292 7760 26298 7772
rect 26418 7760 26424 7772
rect 26476 7760 26482 7812
rect 26881 7803 26939 7809
rect 26881 7769 26893 7803
rect 26927 7800 26939 7803
rect 27062 7800 27068 7812
rect 26927 7772 27068 7800
rect 26927 7769 26939 7772
rect 26881 7763 26939 7769
rect 27062 7760 27068 7772
rect 27120 7760 27126 7812
rect 27540 7744 27568 7831
rect 18984 7704 20668 7732
rect 20717 7735 20775 7741
rect 20717 7701 20729 7735
rect 20763 7732 20775 7735
rect 21174 7732 21180 7744
rect 20763 7704 21180 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 22830 7692 22836 7744
rect 22888 7732 22894 7744
rect 26510 7732 26516 7744
rect 22888 7704 26516 7732
rect 22888 7692 22894 7704
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 27522 7692 27528 7744
rect 27580 7692 27586 7744
rect 27724 7732 27752 7840
rect 27792 7837 27804 7871
rect 27838 7868 27850 7871
rect 28994 7868 29000 7880
rect 27838 7840 29000 7868
rect 27838 7837 27850 7840
rect 27792 7831 27850 7837
rect 28994 7828 29000 7840
rect 29052 7828 29058 7880
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30736 7871 30794 7877
rect 30736 7837 30748 7871
rect 30782 7868 30794 7871
rect 31772 7868 31800 7976
rect 32122 7964 32128 7976
rect 32180 7964 32186 8016
rect 32309 8007 32367 8013
rect 32309 7973 32321 8007
rect 32355 8004 32367 8007
rect 33134 8004 33140 8016
rect 32355 7976 33140 8004
rect 32355 7973 32367 7976
rect 32309 7967 32367 7973
rect 33134 7964 33140 7976
rect 33192 7964 33198 8016
rect 36078 7936 36084 7948
rect 30782 7840 31800 7868
rect 31864 7908 36084 7936
rect 30782 7837 30794 7840
rect 30736 7831 30794 7837
rect 28166 7760 28172 7812
rect 28224 7800 28230 7812
rect 29748 7800 29776 7831
rect 30650 7800 30656 7812
rect 28224 7772 30656 7800
rect 28224 7760 28230 7772
rect 30650 7760 30656 7772
rect 30708 7760 30714 7812
rect 31864 7800 31892 7908
rect 32493 7871 32551 7877
rect 32493 7837 32505 7871
rect 32539 7837 32551 7871
rect 32493 7831 32551 7837
rect 33137 7871 33195 7877
rect 33137 7837 33149 7871
rect 33183 7868 33195 7871
rect 33318 7868 33324 7880
rect 33183 7840 33324 7868
rect 33183 7837 33195 7840
rect 33137 7831 33195 7837
rect 31726 7772 31892 7800
rect 28534 7732 28540 7744
rect 27724 7704 28540 7732
rect 28534 7692 28540 7704
rect 28592 7692 28598 7744
rect 28902 7732 28908 7744
rect 28863 7704 28908 7732
rect 28902 7692 28908 7704
rect 28960 7692 28966 7744
rect 29546 7692 29552 7744
rect 29604 7732 29610 7744
rect 29917 7735 29975 7741
rect 29917 7732 29929 7735
rect 29604 7704 29929 7732
rect 29604 7692 29610 7704
rect 29917 7701 29929 7704
rect 29963 7732 29975 7735
rect 31726 7732 31754 7772
rect 32030 7760 32036 7812
rect 32088 7800 32094 7812
rect 32508 7800 32536 7831
rect 33318 7828 33324 7840
rect 33376 7828 33382 7880
rect 33965 7871 34023 7877
rect 33965 7837 33977 7871
rect 34011 7837 34023 7871
rect 33965 7831 34023 7837
rect 32088 7772 32536 7800
rect 32088 7760 32094 7772
rect 33226 7760 33232 7812
rect 33284 7800 33290 7812
rect 33980 7800 34008 7831
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 35176 7877 35204 7908
rect 36078 7896 36084 7908
rect 36136 7896 36142 7948
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 34848 7840 34897 7868
rect 34848 7828 34854 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 35161 7871 35219 7877
rect 35161 7837 35173 7871
rect 35207 7837 35219 7871
rect 35161 7831 35219 7837
rect 35710 7828 35716 7880
rect 35768 7868 35774 7880
rect 35805 7871 35863 7877
rect 35805 7868 35817 7871
rect 35768 7840 35817 7868
rect 35768 7828 35774 7840
rect 35805 7837 35817 7840
rect 35851 7837 35863 7871
rect 36446 7868 36452 7880
rect 36407 7840 36452 7868
rect 35805 7831 35863 7837
rect 36446 7828 36452 7840
rect 36504 7828 36510 7880
rect 36630 7828 36636 7880
rect 36688 7868 36694 7880
rect 37185 7871 37243 7877
rect 37185 7868 37197 7871
rect 36688 7840 37197 7868
rect 36688 7828 36694 7840
rect 37185 7837 37197 7840
rect 37231 7837 37243 7871
rect 38010 7868 38016 7880
rect 37971 7840 38016 7868
rect 37185 7831 37243 7837
rect 38010 7828 38016 7840
rect 38068 7828 38074 7880
rect 33284 7772 34008 7800
rect 33284 7760 33290 7772
rect 29963 7704 31754 7732
rect 31849 7735 31907 7741
rect 29963 7701 29975 7704
rect 29917 7695 29975 7701
rect 31849 7701 31861 7735
rect 31895 7732 31907 7735
rect 32122 7732 32128 7744
rect 31895 7704 32128 7732
rect 31895 7701 31907 7704
rect 31849 7695 31907 7701
rect 32122 7692 32128 7704
rect 32180 7692 32186 7744
rect 32953 7735 33011 7741
rect 32953 7701 32965 7735
rect 32999 7732 33011 7735
rect 33686 7732 33692 7744
rect 32999 7704 33692 7732
rect 32999 7701 33011 7704
rect 32953 7695 33011 7701
rect 33686 7692 33692 7704
rect 33744 7692 33750 7744
rect 34698 7732 34704 7744
rect 34659 7704 34704 7732
rect 34698 7692 34704 7704
rect 34756 7692 34762 7744
rect 35069 7735 35127 7741
rect 35069 7701 35081 7735
rect 35115 7732 35127 7735
rect 35434 7732 35440 7744
rect 35115 7704 35440 7732
rect 35115 7701 35127 7704
rect 35069 7695 35127 7701
rect 35434 7692 35440 7704
rect 35492 7692 35498 7744
rect 35618 7732 35624 7744
rect 35579 7704 35624 7732
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 36262 7732 36268 7744
rect 36223 7704 36268 7732
rect 36262 7692 36268 7704
rect 36320 7692 36326 7744
rect 37001 7735 37059 7741
rect 37001 7701 37013 7735
rect 37047 7732 37059 7735
rect 37642 7732 37648 7744
rect 37047 7704 37648 7732
rect 37047 7701 37059 7704
rect 37001 7695 37059 7701
rect 37642 7692 37648 7704
rect 37700 7692 37706 7744
rect 37826 7732 37832 7744
rect 37787 7704 37832 7732
rect 37826 7692 37832 7704
rect 37884 7692 37890 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 3694 7528 3700 7540
rect 3655 7500 3700 7528
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 10226 7528 10232 7540
rect 6880 7500 10232 7528
rect 6880 7488 6886 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 11606 7528 11612 7540
rect 10336 7500 11612 7528
rect 6733 7463 6791 7469
rect 6733 7460 6745 7463
rect 6196 7432 6745 7460
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 992 7364 1593 7392
rect 992 7352 998 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 2593 7355 2651 7361
rect 2608 7324 2636 7355
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 4430 7392 4436 7404
rect 3927 7364 4436 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5350 7392 5356 7404
rect 5215 7364 5356 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 3970 7324 3976 7336
rect 2608 7296 3976 7324
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4540 7324 4568 7355
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6196 7392 6224 7432
rect 6733 7429 6745 7432
rect 6779 7429 6791 7463
rect 6733 7423 6791 7429
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 7438 7463 7496 7469
rect 7438 7460 7450 7463
rect 6972 7432 7450 7460
rect 6972 7420 6978 7432
rect 7438 7429 7450 7432
rect 7484 7429 7496 7463
rect 7438 7423 7496 7429
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 10336 7460 10364 7500
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 14274 7528 14280 7540
rect 11992 7500 14280 7528
rect 7892 7432 10364 7460
rect 10965 7463 11023 7469
rect 7892 7420 7898 7432
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11992 7460 12020 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 14734 7528 14740 7540
rect 14608 7500 14740 7528
rect 14608 7488 14614 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15194 7528 15200 7540
rect 15155 7500 15200 7528
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 23014 7528 23020 7540
rect 22572 7500 23020 7528
rect 11011 7432 12020 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12774 7463 12832 7469
rect 12774 7460 12786 7463
rect 12124 7432 12786 7460
rect 12124 7420 12130 7432
rect 12774 7429 12786 7432
rect 12820 7429 12832 7463
rect 15654 7460 15660 7472
rect 12774 7423 12832 7429
rect 14660 7432 15660 7460
rect 6362 7392 6368 7404
rect 5859 7364 6224 7392
rect 6323 7364 6368 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6549 7396 6607 7401
rect 6549 7395 6684 7396
rect 6549 7361 6561 7395
rect 6595 7392 6684 7395
rect 7006 7392 7012 7404
rect 6595 7368 7012 7392
rect 6595 7361 6607 7368
rect 6656 7364 7012 7368
rect 6549 7355 6607 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8536 7364 9045 7392
rect 8536 7352 8542 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9033 7355 9091 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 10134 7392 10140 7404
rect 10095 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11054 7392 11060 7404
rect 10827 7364 11060 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11701 7395 11759 7401
rect 11204 7364 11652 7392
rect 11204 7352 11210 7364
rect 6822 7324 6828 7336
rect 4540 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 6972 7296 7205 7324
rect 6972 7284 6978 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 7193 7287 7251 7293
rect 8220 7296 9137 7324
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 5166 7256 5172 7268
rect 2455 7228 5172 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 5592 7228 5641 7256
rect 5592 7216 5598 7228
rect 5629 7225 5641 7228
rect 5675 7225 5687 7259
rect 5629 7219 5687 7225
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 1762 7188 1768 7200
rect 1443 7160 1768 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4890 7188 4896 7200
rect 4387 7160 4896 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 4985 7191 5043 7197
rect 4985 7157 4997 7191
rect 5031 7188 5043 7191
rect 6362 7188 6368 7200
rect 5031 7160 6368 7188
rect 5031 7157 5043 7160
rect 4985 7151 5043 7157
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8220 7188 8248 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9784 7324 9812 7352
rect 10042 7324 10048 7336
rect 9784 7296 10048 7324
rect 9125 7287 9183 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10594 7324 10600 7336
rect 10507 7296 10600 7324
rect 10594 7284 10600 7296
rect 10652 7324 10658 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 10652 7296 11529 7324
rect 10652 7284 10658 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11624 7324 11652 7364
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12250 7392 12256 7404
rect 11747 7364 12256 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 13998 7392 14004 7404
rect 12406 7364 14004 7392
rect 12158 7324 12164 7336
rect 11624 7296 12164 7324
rect 11517 7287 11575 7293
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8352 7228 10180 7256
rect 8352 7216 8358 7228
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8168 7160 8585 7188
rect 8168 7148 8174 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 9030 7188 9036 7200
rect 8991 7160 9036 7188
rect 8573 7151 8631 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 9364 7160 9505 7188
rect 9364 7148 9370 7160
rect 9493 7157 9505 7160
rect 9539 7157 9551 7191
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9493 7151 9551 7157
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10152 7188 10180 7228
rect 10226 7216 10232 7268
rect 10284 7256 10290 7268
rect 12406 7256 12434 7364
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14660 7401 14688 7432
rect 15212 7404 15240 7432
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 17129 7463 17187 7469
rect 17129 7460 17141 7463
rect 16632 7432 17141 7460
rect 16632 7420 16638 7432
rect 17129 7429 17141 7432
rect 17175 7460 17187 7463
rect 17586 7460 17592 7472
rect 17175 7432 17592 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 17957 7463 18015 7469
rect 17957 7429 17969 7463
rect 18003 7460 18015 7463
rect 18414 7460 18420 7472
rect 18003 7432 18420 7460
rect 18003 7429 18015 7432
rect 17957 7423 18015 7429
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 22094 7460 22100 7472
rect 19904 7432 22100 7460
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7361 14703 7395
rect 14826 7392 14832 7404
rect 14787 7364 14832 7392
rect 14645 7355 14703 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12584 7296 12629 7324
rect 12584 7284 12590 7296
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14936 7324 14964 7355
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 15068 7364 15113 7392
rect 15068 7352 15074 7364
rect 15194 7352 15200 7404
rect 15252 7352 15258 7404
rect 15838 7392 15844 7404
rect 15799 7364 15844 7392
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17276 7364 17785 7392
rect 17276 7352 17282 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18187 7364 18797 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18785 7361 18797 7364
rect 18831 7361 18843 7395
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 18785 7355 18843 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19904 7401 19932 7432
rect 22094 7420 22100 7432
rect 22152 7460 22158 7472
rect 22370 7460 22376 7472
rect 22152 7432 22376 7460
rect 22152 7420 22158 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 20156 7395 20214 7401
rect 20156 7361 20168 7395
rect 20202 7392 20214 7395
rect 20530 7392 20536 7404
rect 20202 7364 20536 7392
rect 20202 7361 20214 7364
rect 20156 7355 20214 7361
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22572 7392 22600 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 28537 7531 28595 7537
rect 28537 7528 28549 7531
rect 24728 7500 28549 7528
rect 24728 7488 24734 7500
rect 28537 7497 28549 7500
rect 28583 7497 28595 7531
rect 28537 7491 28595 7497
rect 28626 7488 28632 7540
rect 28684 7528 28690 7540
rect 31389 7531 31447 7537
rect 28684 7500 31340 7528
rect 28684 7488 28690 7500
rect 23845 7463 23903 7469
rect 23845 7429 23857 7463
rect 23891 7460 23903 7463
rect 24578 7460 24584 7472
rect 23891 7432 24584 7460
rect 23891 7429 23903 7432
rect 23845 7423 23903 7429
rect 24578 7420 24584 7432
rect 24636 7420 24642 7472
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 27614 7460 27620 7472
rect 26936 7432 27476 7460
rect 27575 7432 27620 7460
rect 26936 7420 26942 7432
rect 22235 7364 22600 7392
rect 23109 7396 23167 7401
rect 23109 7395 23244 7396
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 23109 7361 23121 7395
rect 23155 7392 23244 7395
rect 23934 7392 23940 7404
rect 23155 7368 23940 7392
rect 23155 7361 23167 7368
rect 23216 7364 23940 7368
rect 23109 7355 23167 7361
rect 23934 7352 23940 7364
rect 23992 7352 23998 7404
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24084 7364 24685 7392
rect 24084 7352 24090 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24762 7352 24768 7404
rect 24820 7392 24826 7404
rect 25041 7395 25099 7401
rect 24820 7364 24865 7392
rect 24820 7352 24826 7364
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25590 7392 25596 7404
rect 25087 7364 25596 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 25685 7395 25743 7401
rect 25685 7361 25697 7395
rect 25731 7392 25743 7395
rect 26142 7392 26148 7404
rect 25731 7364 26148 7392
rect 25731 7361 25743 7364
rect 25685 7355 25743 7361
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 26418 7392 26424 7404
rect 26379 7364 26424 7392
rect 26418 7352 26424 7364
rect 26476 7352 26482 7404
rect 26510 7352 26516 7404
rect 26568 7392 26574 7404
rect 27448 7401 27476 7432
rect 27614 7420 27620 7432
rect 27672 7420 27678 7472
rect 28902 7460 28908 7472
rect 27816 7432 28908 7460
rect 27816 7401 27844 7432
rect 28902 7420 28908 7432
rect 28960 7420 28966 7472
rect 29448 7463 29506 7469
rect 29448 7429 29460 7463
rect 29494 7460 29506 7463
rect 30282 7460 30288 7472
rect 29494 7432 30288 7460
rect 29494 7429 29506 7432
rect 29448 7423 29506 7429
rect 30282 7420 30288 7432
rect 30340 7420 30346 7472
rect 31021 7463 31079 7469
rect 31021 7429 31033 7463
rect 31067 7429 31079 7463
rect 31021 7423 31079 7429
rect 27249 7395 27307 7401
rect 27249 7392 27261 7395
rect 26568 7364 27261 7392
rect 26568 7352 26574 7364
rect 27249 7361 27261 7364
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7392 27951 7395
rect 28166 7392 28172 7404
rect 27939 7364 28172 7392
rect 27939 7361 27951 7364
rect 27893 7355 27951 7361
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7361 28779 7395
rect 29178 7392 29184 7404
rect 29139 7364 29184 7392
rect 28721 7355 28779 7361
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 14424 7296 14964 7324
rect 15212 7296 15669 7324
rect 14424 7284 14430 7296
rect 14826 7256 14832 7268
rect 10284 7228 12434 7256
rect 13740 7228 14832 7256
rect 10284 7216 10290 7228
rect 12066 7188 12072 7200
rect 10152 7160 12072 7188
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13740 7188 13768 7228
rect 14826 7216 14832 7228
rect 14884 7256 14890 7268
rect 15102 7256 15108 7268
rect 14884 7228 15108 7256
rect 14884 7216 14890 7228
rect 15102 7216 15108 7228
rect 15160 7216 15166 7268
rect 13906 7188 13912 7200
rect 13320 7160 13768 7188
rect 13867 7160 13912 7188
rect 13320 7148 13326 7160
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 15212 7188 15240 7296
rect 15657 7293 15669 7296
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7324 22431 7327
rect 28736 7324 28764 7355
rect 29178 7352 29184 7364
rect 29236 7352 29242 7404
rect 31036 7392 31064 7423
rect 31110 7420 31116 7472
rect 31168 7460 31174 7472
rect 31221 7463 31279 7469
rect 31221 7460 31233 7463
rect 31168 7432 31233 7460
rect 31168 7420 31174 7432
rect 31221 7429 31233 7432
rect 31267 7429 31279 7463
rect 31312 7460 31340 7500
rect 31389 7497 31401 7531
rect 31435 7528 31447 7531
rect 32306 7528 32312 7540
rect 31435 7500 32312 7528
rect 31435 7497 31447 7500
rect 31389 7491 31447 7497
rect 32306 7488 32312 7500
rect 32364 7488 32370 7540
rect 32392 7463 32450 7469
rect 31312 7432 32352 7460
rect 31221 7423 31279 7429
rect 32324 7392 32352 7432
rect 32392 7429 32404 7463
rect 32438 7460 32450 7463
rect 32766 7460 32772 7472
rect 32438 7432 32772 7460
rect 32438 7429 32450 7432
rect 32392 7423 32450 7429
rect 32766 7420 32772 7432
rect 32824 7420 32830 7472
rect 34232 7463 34290 7469
rect 34232 7429 34244 7463
rect 34278 7460 34290 7463
rect 34698 7460 34704 7472
rect 34278 7432 34704 7460
rect 34278 7429 34290 7432
rect 34232 7423 34290 7429
rect 34698 7420 34704 7432
rect 34756 7420 34762 7472
rect 36078 7420 36084 7472
rect 36136 7460 36142 7472
rect 36136 7432 36308 7460
rect 36136 7420 36142 7432
rect 33594 7392 33600 7404
rect 31036 7364 31800 7392
rect 32324 7364 33600 7392
rect 22419 7296 28764 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 19886 7256 19892 7268
rect 17236 7228 19892 7256
rect 14240 7160 15240 7188
rect 14240 7148 14246 7160
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 17236 7197 17264 7228
rect 19886 7216 19892 7228
rect 19944 7216 19950 7268
rect 22278 7216 22284 7268
rect 22336 7256 22342 7268
rect 23382 7256 23388 7268
rect 22336 7228 23388 7256
rect 22336 7216 22342 7228
rect 23382 7216 23388 7228
rect 23440 7256 23446 7268
rect 24949 7259 25007 7265
rect 23440 7228 24900 7256
rect 23440 7216 23446 7228
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 16540 7160 17233 7188
rect 16540 7148 16546 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 18598 7188 18604 7200
rect 18559 7160 18604 7188
rect 17221 7151 17279 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 19245 7191 19303 7197
rect 19245 7157 19257 7191
rect 19291 7188 19303 7191
rect 19334 7188 19340 7200
rect 19291 7160 19340 7188
rect 19291 7157 19303 7160
rect 19245 7151 19303 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 22830 7148 22836 7200
rect 22888 7188 22894 7200
rect 22925 7191 22983 7197
rect 22925 7188 22937 7191
rect 22888 7160 22937 7188
rect 22888 7148 22894 7160
rect 22925 7157 22937 7160
rect 22971 7157 22983 7191
rect 22925 7151 22983 7157
rect 23937 7191 23995 7197
rect 23937 7157 23949 7191
rect 23983 7188 23995 7191
rect 24302 7188 24308 7200
rect 23983 7160 24308 7188
rect 23983 7157 23995 7160
rect 23937 7151 23995 7157
rect 24302 7148 24308 7160
rect 24360 7148 24366 7200
rect 24394 7148 24400 7200
rect 24452 7188 24458 7200
rect 24489 7191 24547 7197
rect 24489 7188 24501 7191
rect 24452 7160 24501 7188
rect 24452 7148 24458 7160
rect 24489 7157 24501 7160
rect 24535 7157 24547 7191
rect 24872 7188 24900 7228
rect 24949 7225 24961 7259
rect 24995 7256 25007 7259
rect 25130 7256 25136 7268
rect 24995 7228 25136 7256
rect 24995 7225 25007 7228
rect 24949 7219 25007 7225
rect 25130 7216 25136 7228
rect 25188 7216 25194 7268
rect 26237 7259 26295 7265
rect 25332 7228 26188 7256
rect 25332 7188 25360 7228
rect 25498 7188 25504 7200
rect 24872 7160 25360 7188
rect 25459 7160 25504 7188
rect 24489 7151 24547 7157
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 26160 7188 26188 7228
rect 26237 7225 26249 7259
rect 26283 7256 26295 7259
rect 28350 7256 28356 7268
rect 26283 7228 28356 7256
rect 26283 7225 26295 7228
rect 26237 7219 26295 7225
rect 28350 7216 28356 7228
rect 28408 7216 28414 7268
rect 29546 7188 29552 7200
rect 26160 7160 29552 7188
rect 29546 7148 29552 7160
rect 29604 7148 29610 7200
rect 29822 7148 29828 7200
rect 29880 7188 29886 7200
rect 30561 7191 30619 7197
rect 30561 7188 30573 7191
rect 29880 7160 30573 7188
rect 29880 7148 29886 7160
rect 30561 7157 30573 7160
rect 30607 7157 30619 7191
rect 31202 7188 31208 7200
rect 31163 7160 31208 7188
rect 30561 7151 30619 7157
rect 31202 7148 31208 7160
rect 31260 7148 31266 7200
rect 31772 7188 31800 7364
rect 33594 7352 33600 7364
rect 33652 7352 33658 7404
rect 34790 7352 34796 7404
rect 34848 7392 34854 7404
rect 35989 7395 36047 7401
rect 35989 7392 36001 7395
rect 34848 7364 36001 7392
rect 34848 7352 34854 7364
rect 35989 7361 36001 7364
rect 36035 7361 36047 7395
rect 36170 7392 36176 7404
rect 36131 7364 36176 7392
rect 35989 7355 36047 7361
rect 36170 7352 36176 7364
rect 36228 7352 36234 7404
rect 36280 7401 36308 7432
rect 36265 7395 36323 7401
rect 36265 7361 36277 7395
rect 36311 7392 36323 7395
rect 36814 7392 36820 7404
rect 36311 7364 36820 7392
rect 36311 7361 36323 7364
rect 36265 7355 36323 7361
rect 36814 7352 36820 7364
rect 36872 7352 36878 7404
rect 36906 7352 36912 7404
rect 36964 7392 36970 7404
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 36964 7364 37473 7392
rect 36964 7352 36970 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 38102 7392 38108 7404
rect 38063 7364 38108 7392
rect 37461 7355 37519 7361
rect 38102 7352 38108 7364
rect 38160 7352 38166 7404
rect 31938 7284 31944 7336
rect 31996 7324 32002 7336
rect 32125 7327 32183 7333
rect 32125 7324 32137 7327
rect 31996 7296 32137 7324
rect 31996 7284 32002 7296
rect 32125 7293 32137 7296
rect 32171 7293 32183 7327
rect 33962 7324 33968 7336
rect 33923 7296 33968 7324
rect 32125 7287 32183 7293
rect 33962 7284 33968 7296
rect 34020 7284 34026 7336
rect 36722 7216 36728 7268
rect 36780 7256 36786 7268
rect 37921 7259 37979 7265
rect 37921 7256 37933 7259
rect 36780 7228 37933 7256
rect 36780 7216 36786 7228
rect 37921 7225 37933 7228
rect 37967 7225 37979 7259
rect 37921 7219 37979 7225
rect 32122 7188 32128 7200
rect 31772 7160 32128 7188
rect 32122 7148 32128 7160
rect 32180 7148 32186 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 33505 7191 33563 7197
rect 33505 7188 33517 7191
rect 32456 7160 33517 7188
rect 32456 7148 32462 7160
rect 33505 7157 33517 7160
rect 33551 7157 33563 7191
rect 33505 7151 33563 7157
rect 35345 7191 35403 7197
rect 35345 7157 35357 7191
rect 35391 7188 35403 7191
rect 35434 7188 35440 7200
rect 35391 7160 35440 7188
rect 35391 7157 35403 7160
rect 35345 7151 35403 7157
rect 35434 7148 35440 7160
rect 35492 7148 35498 7200
rect 35802 7188 35808 7200
rect 35763 7160 35808 7188
rect 35802 7148 35808 7160
rect 35860 7148 35866 7200
rect 37274 7188 37280 7200
rect 37235 7160 37280 7188
rect 37274 7148 37280 7160
rect 37332 7148 37338 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 2958 6984 2964 6996
rect 2919 6956 2964 6984
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3108 6956 7052 6984
rect 3108 6944 3114 6956
rect 1673 6919 1731 6925
rect 1673 6885 1685 6919
rect 1719 6914 1731 6919
rect 4522 6916 4528 6928
rect 1719 6886 1753 6914
rect 2792 6888 4528 6916
rect 1719 6885 1731 6886
rect 1673 6879 1731 6885
rect 1688 6848 1716 6879
rect 2792 6848 2820 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 7024 6916 7052 6956
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7156 6956 7941 6984
rect 7156 6944 7162 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 8846 6944 8852 6996
rect 8904 6984 8910 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 8904 6956 9137 6984
rect 8904 6944 8910 6956
rect 9125 6953 9137 6956
rect 9171 6953 9183 6987
rect 9125 6947 9183 6953
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10594 6984 10600 6996
rect 9732 6956 10600 6984
rect 9732 6944 9738 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 10778 6984 10784 6996
rect 10739 6956 10784 6984
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 12342 6984 12348 6996
rect 12303 6956 12348 6984
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13170 6984 13176 6996
rect 12492 6956 13176 6984
rect 12492 6944 12498 6956
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 14366 6984 14372 6996
rect 14327 6956 14372 6984
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 15988 6956 19334 6984
rect 15988 6944 15994 6956
rect 13446 6916 13452 6928
rect 4764 6888 4809 6916
rect 7024 6888 13452 6916
rect 4764 6876 4770 6888
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 13722 6876 13728 6928
rect 13780 6916 13786 6928
rect 18325 6919 18383 6925
rect 13780 6888 14044 6916
rect 13780 6876 13786 6888
rect 1688 6820 2820 6848
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 5442 6848 5448 6860
rect 3936 6820 5448 6848
rect 3936 6808 3942 6820
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5500 6820 5549 6848
rect 5500 6808 5506 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 7248 6820 9229 6848
rect 7248 6808 7254 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9950 6848 9956 6860
rect 9732 6820 9956 6848
rect 9732 6808 9738 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10744 6820 10793 6848
rect 10744 6808 10750 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12618 6848 12624 6860
rect 12299 6820 12624 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 13906 6848 13912 6860
rect 13004 6820 13912 6848
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 2406 6780 2412 6792
rect 1903 6752 2412 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2774 6780 2780 6792
rect 2547 6752 2780 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3234 6780 3240 6792
rect 3191 6752 3240 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4798 6780 4804 6792
rect 4295 6752 4804 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6749 4951 6783
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 4893 6743 4951 6749
rect 7024 6752 7389 6780
rect 4908 6656 4936 6743
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 5782 6715 5840 6721
rect 5782 6712 5794 6715
rect 5592 6684 5794 6712
rect 5592 6672 5598 6684
rect 5782 6681 5794 6684
rect 5828 6681 5840 6715
rect 5782 6675 5840 6681
rect 5902 6672 5908 6724
rect 5960 6712 5966 6724
rect 6546 6712 6552 6724
rect 5960 6684 6552 6712
rect 5960 6672 5966 6684
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 7024 6656 7052 6752
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7377 6743 7435 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9306 6780 9312 6792
rect 9171 6752 9312 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9582 6780 9588 6792
rect 9447 6752 9588 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11238 6780 11244 6792
rect 11011 6752 11244 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 12894 6780 12900 6792
rect 12391 6752 12900 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13004 6789 13032 6820
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14016 6848 14044 6888
rect 18325 6885 18337 6919
rect 18371 6885 18383 6919
rect 19306 6916 19334 6956
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 19484 6956 19901 6984
rect 19484 6944 19490 6956
rect 19889 6953 19901 6956
rect 19935 6953 19947 6987
rect 19889 6947 19947 6953
rect 20809 6987 20867 6993
rect 20809 6953 20821 6987
rect 20855 6984 20867 6987
rect 22646 6984 22652 6996
rect 20855 6956 22652 6984
rect 20855 6953 20867 6956
rect 20809 6947 20867 6953
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 27890 6944 27896 6996
rect 27948 6984 27954 6996
rect 31570 6984 31576 6996
rect 27948 6956 31576 6984
rect 27948 6944 27954 6956
rect 31570 6944 31576 6956
rect 31628 6944 31634 6996
rect 23106 6916 23112 6928
rect 19306 6888 23112 6916
rect 18325 6879 18383 6885
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14016 6820 14197 6848
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 18340 6848 18368 6879
rect 20990 6848 20996 6860
rect 18340 6820 20996 6848
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 13136 6752 13277 6780
rect 13136 6740 13142 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13630 6780 13636 6792
rect 13403 6752 13636 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13924 6780 13952 6808
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13924 6752 14381 6780
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 15059 6752 16957 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 16945 6749 16957 6752
rect 16991 6780 17003 6783
rect 18046 6780 18052 6792
rect 16991 6752 18052 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 7282 6672 7288 6724
rect 7340 6712 7346 6724
rect 7561 6715 7619 6721
rect 7561 6712 7573 6715
rect 7340 6684 7573 6712
rect 7340 6672 7346 6684
rect 7561 6681 7573 6684
rect 7607 6681 7619 6715
rect 7561 6675 7619 6681
rect 7653 6715 7711 6721
rect 7653 6681 7665 6715
rect 7699 6712 7711 6715
rect 7834 6712 7840 6724
rect 7699 6684 7840 6712
rect 7699 6681 7711 6684
rect 7653 6675 7711 6681
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4890 6604 4896 6656
rect 4948 6604 4954 6656
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 6822 6644 6828 6656
rect 5040 6616 6828 6644
rect 5040 6604 5046 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7006 6644 7012 6656
rect 6963 6616 7012 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7576 6644 7604 6675
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 10318 6712 10324 6724
rect 8720 6684 10324 6712
rect 8720 6672 8726 6684
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10502 6672 10508 6724
rect 10560 6712 10566 6724
rect 10689 6715 10747 6721
rect 10689 6712 10701 6715
rect 10560 6684 10701 6712
rect 10560 6672 10566 6684
rect 10689 6681 10701 6684
rect 10735 6681 10747 6715
rect 10689 6675 10747 6681
rect 10980 6684 12020 6712
rect 7926 6644 7932 6656
rect 7576 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 10980 6644 11008 6684
rect 11146 6644 11152 6656
rect 9631 6616 11008 6644
rect 11107 6616 11152 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11992 6644 12020 6684
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12802 6712 12808 6724
rect 12124 6684 12169 6712
rect 12406 6684 12808 6712
rect 12124 6672 12130 6684
rect 12406 6644 12434 6684
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6681 13231 6715
rect 14090 6712 14096 6724
rect 14051 6684 14096 6712
rect 13173 6675 13231 6681
rect 11992 6616 12434 6644
rect 12529 6647 12587 6653
rect 12529 6613 12541 6647
rect 12575 6644 12587 6647
rect 13078 6644 13084 6656
rect 12575 6616 13084 6644
rect 12575 6613 12587 6616
rect 12529 6607 12587 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13188 6644 13216 6675
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 15028 6712 15056 6743
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 14240 6684 15056 6712
rect 15280 6715 15338 6721
rect 14240 6672 14246 6684
rect 15280 6681 15292 6715
rect 15326 6712 15338 6715
rect 15746 6712 15752 6724
rect 15326 6684 15752 6712
rect 15326 6681 15338 6684
rect 15280 6675 15338 6681
rect 15746 6672 15752 6684
rect 15804 6672 15810 6724
rect 15930 6672 15936 6724
rect 15988 6712 15994 6724
rect 17190 6715 17248 6721
rect 17190 6712 17202 6715
rect 15988 6684 17202 6712
rect 15988 6672 15994 6684
rect 17190 6681 17202 6684
rect 17236 6681 17248 6715
rect 17190 6675 17248 6681
rect 17862 6672 17868 6724
rect 17920 6712 17926 6724
rect 18340 6712 18368 6820
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 19978 6780 19984 6792
rect 19567 6752 19984 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 21560 6789 21588 6888
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 23201 6919 23259 6925
rect 23201 6885 23213 6919
rect 23247 6916 23259 6919
rect 23290 6916 23296 6928
rect 23247 6888 23296 6916
rect 23247 6885 23259 6888
rect 23201 6879 23259 6885
rect 23290 6876 23296 6888
rect 23348 6876 23354 6928
rect 25590 6876 25596 6928
rect 25648 6916 25654 6928
rect 25869 6919 25927 6925
rect 25869 6916 25881 6919
rect 25648 6888 25881 6916
rect 25648 6876 25654 6888
rect 25869 6885 25881 6888
rect 25915 6885 25927 6919
rect 25869 6879 25927 6885
rect 26804 6888 28028 6916
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22152 6820 22784 6848
rect 22152 6808 22158 6820
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6780 21787 6783
rect 22002 6780 22008 6792
rect 21775 6752 22008 6780
rect 21775 6749 21787 6752
rect 21729 6743 21787 6749
rect 22002 6740 22008 6752
rect 22060 6740 22066 6792
rect 22278 6740 22284 6792
rect 22336 6780 22342 6792
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 22336 6752 22385 6780
rect 22336 6740 22342 6752
rect 22373 6749 22385 6752
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 22646 6780 22652 6792
rect 22603 6752 22652 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 22756 6780 22784 6820
rect 26234 6808 26240 6860
rect 26292 6848 26298 6860
rect 26510 6848 26516 6860
rect 26292 6820 26516 6848
rect 26292 6808 26298 6820
rect 26510 6808 26516 6820
rect 26568 6848 26574 6860
rect 26605 6851 26663 6857
rect 26605 6848 26617 6851
rect 26568 6820 26617 6848
rect 26568 6808 26574 6820
rect 26605 6817 26617 6820
rect 26651 6817 26663 6851
rect 26804 6848 26832 6888
rect 26605 6811 26663 6817
rect 26712 6820 26832 6848
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22756 6752 23029 6780
rect 23017 6749 23029 6752
rect 23063 6780 23075 6783
rect 23566 6780 23572 6792
rect 23063 6752 23572 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 24302 6740 24308 6792
rect 24360 6780 24366 6792
rect 24489 6783 24547 6789
rect 24489 6780 24501 6783
rect 24360 6752 24501 6780
rect 24360 6740 24366 6752
rect 24489 6749 24501 6752
rect 24535 6749 24547 6783
rect 24489 6743 24547 6749
rect 24756 6783 24814 6789
rect 24756 6749 24768 6783
rect 24802 6780 24814 6783
rect 26712 6780 26740 6820
rect 26878 6808 26884 6860
rect 26936 6848 26942 6860
rect 26936 6820 27752 6848
rect 26936 6808 26942 6820
rect 24802 6752 26740 6780
rect 26789 6783 26847 6789
rect 24802 6749 24814 6752
rect 24756 6743 24814 6749
rect 26789 6749 26801 6783
rect 26835 6780 26847 6783
rect 26896 6780 26924 6808
rect 26835 6752 26924 6780
rect 26993 6761 27051 6767
rect 26835 6749 26847 6752
rect 26789 6743 26847 6749
rect 26993 6727 27005 6761
rect 27039 6758 27051 6761
rect 27039 6727 27052 6758
rect 27430 6740 27436 6792
rect 27488 6780 27494 6792
rect 27724 6789 27752 6820
rect 27798 6808 27804 6860
rect 27856 6848 27862 6860
rect 28000 6848 28028 6888
rect 28810 6848 28816 6860
rect 27856 6820 27901 6848
rect 28000 6820 28816 6848
rect 27856 6808 27862 6820
rect 28810 6808 28816 6820
rect 28868 6808 28874 6860
rect 29178 6808 29184 6860
rect 29236 6848 29242 6860
rect 29549 6851 29607 6857
rect 29549 6848 29561 6851
rect 29236 6820 29561 6848
rect 29236 6808 29242 6820
rect 29549 6817 29561 6820
rect 29595 6817 29607 6851
rect 29549 6811 29607 6817
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 30616 6820 32076 6848
rect 30616 6808 30622 6820
rect 27525 6783 27583 6789
rect 27525 6780 27537 6783
rect 27488 6752 27537 6780
rect 27488 6740 27494 6752
rect 27525 6749 27537 6752
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6749 27767 6783
rect 27709 6743 27767 6749
rect 27898 6783 27956 6789
rect 27898 6749 27910 6783
rect 27944 6780 27956 6783
rect 28166 6780 28172 6792
rect 27944 6752 28172 6780
rect 27944 6749 27972 6752
rect 27898 6743 27972 6749
rect 17920 6684 18368 6712
rect 17920 6672 17926 6684
rect 18414 6672 18420 6724
rect 18472 6712 18478 6724
rect 19705 6715 19763 6721
rect 19705 6712 19717 6715
rect 18472 6684 19717 6712
rect 18472 6672 18478 6684
rect 19705 6681 19717 6684
rect 19751 6712 19763 6715
rect 20530 6712 20536 6724
rect 19751 6684 20536 6712
rect 19751 6681 19763 6684
rect 19705 6675 19763 6681
rect 20530 6672 20536 6684
rect 20588 6672 20594 6724
rect 20714 6712 20720 6724
rect 20627 6684 20720 6712
rect 20714 6672 20720 6684
rect 20772 6712 20778 6724
rect 21821 6715 21879 6721
rect 21821 6712 21833 6715
rect 20772 6684 21833 6712
rect 20772 6672 20778 6684
rect 21821 6681 21833 6684
rect 21867 6681 21879 6715
rect 21821 6675 21879 6681
rect 21913 6715 21971 6721
rect 21913 6681 21925 6715
rect 21959 6712 21971 6715
rect 22922 6712 22928 6724
rect 21959 6684 22928 6712
rect 21959 6681 21971 6684
rect 21913 6675 21971 6681
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 26605 6715 26663 6721
rect 26605 6681 26617 6715
rect 26651 6681 26663 6715
rect 26878 6712 26884 6724
rect 26839 6684 26884 6712
rect 26605 6675 26663 6681
rect 13262 6644 13268 6656
rect 13188 6616 13268 6644
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 13538 6644 13544 6656
rect 13499 6616 13544 6644
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 16264 6616 16405 6644
rect 16264 6604 16270 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 20346 6644 20352 6656
rect 16724 6616 20352 6644
rect 16724 6604 16730 6616
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 22554 6644 22560 6656
rect 22515 6616 22560 6644
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 26620 6644 26648 6675
rect 26878 6672 26884 6684
rect 26936 6672 26942 6724
rect 26993 6721 27052 6727
rect 27024 6712 27052 6721
rect 27024 6684 27108 6712
rect 26970 6644 26976 6656
rect 26620 6616 26976 6644
rect 26970 6604 26976 6616
rect 27028 6604 27034 6656
rect 27080 6644 27108 6684
rect 27798 6672 27804 6724
rect 27856 6712 27862 6724
rect 27856 6684 27901 6712
rect 27856 6672 27862 6684
rect 27944 6644 27972 6743
rect 28166 6740 28172 6752
rect 28224 6740 28230 6792
rect 28534 6780 28540 6792
rect 28495 6752 28540 6780
rect 28534 6740 28540 6752
rect 28592 6740 28598 6792
rect 29816 6783 29874 6789
rect 29816 6749 29828 6783
rect 29862 6780 29874 6783
rect 30190 6780 30196 6792
rect 29862 6752 30196 6780
rect 29862 6749 29874 6752
rect 29816 6743 29874 6749
rect 30190 6740 30196 6752
rect 30248 6740 30254 6792
rect 31938 6780 31944 6792
rect 31851 6752 31944 6780
rect 31938 6740 31944 6752
rect 31996 6740 32002 6792
rect 32048 6780 32076 6820
rect 33873 6783 33931 6789
rect 33873 6780 33885 6783
rect 32048 6752 33885 6780
rect 33873 6749 33885 6752
rect 33919 6749 33931 6783
rect 33873 6743 33931 6749
rect 34057 6783 34115 6789
rect 34057 6749 34069 6783
rect 34103 6780 34115 6783
rect 34698 6780 34704 6792
rect 34103 6752 34704 6780
rect 34103 6749 34115 6752
rect 34057 6743 34115 6749
rect 28721 6715 28779 6721
rect 28721 6681 28733 6715
rect 28767 6712 28779 6715
rect 30742 6712 30748 6724
rect 28767 6684 30748 6712
rect 28767 6681 28779 6684
rect 28721 6675 28779 6681
rect 30742 6672 30748 6684
rect 30800 6712 30806 6724
rect 31662 6712 31668 6724
rect 30800 6684 31668 6712
rect 30800 6672 30806 6684
rect 31662 6672 31668 6684
rect 31720 6672 31726 6724
rect 27080 6616 27972 6644
rect 29270 6604 29276 6656
rect 29328 6644 29334 6656
rect 30929 6647 30987 6653
rect 30929 6644 30941 6647
rect 29328 6616 30941 6644
rect 29328 6604 29334 6616
rect 30929 6613 30941 6616
rect 30975 6613 30987 6647
rect 30929 6607 30987 6613
rect 31294 6604 31300 6656
rect 31352 6644 31358 6656
rect 31846 6644 31852 6656
rect 31352 6616 31852 6644
rect 31352 6604 31358 6616
rect 31846 6604 31852 6616
rect 31904 6604 31910 6656
rect 31956 6644 31984 6740
rect 32214 6721 32220 6724
rect 32208 6712 32220 6721
rect 32175 6684 32220 6712
rect 32208 6675 32220 6684
rect 32214 6672 32220 6675
rect 32272 6672 32278 6724
rect 33962 6712 33968 6724
rect 32324 6684 33968 6712
rect 32324 6644 32352 6684
rect 33962 6672 33968 6684
rect 34020 6712 34026 6724
rect 34072 6712 34100 6743
rect 34698 6740 34704 6752
rect 34756 6740 34762 6792
rect 36725 6783 36783 6789
rect 36725 6780 36737 6783
rect 34900 6752 36737 6780
rect 34020 6684 34100 6712
rect 34020 6672 34026 6684
rect 34790 6672 34796 6724
rect 34848 6712 34854 6724
rect 34900 6712 34928 6752
rect 36725 6749 36737 6752
rect 36771 6749 36783 6783
rect 36725 6743 36783 6749
rect 36814 6740 36820 6792
rect 36872 6780 36878 6792
rect 37001 6783 37059 6789
rect 37001 6780 37013 6783
rect 36872 6752 37013 6780
rect 36872 6740 36878 6752
rect 37001 6749 37013 6752
rect 37047 6749 37059 6783
rect 37001 6743 37059 6749
rect 37182 6740 37188 6792
rect 37240 6780 37246 6792
rect 37645 6783 37703 6789
rect 37645 6780 37657 6783
rect 37240 6752 37657 6780
rect 37240 6740 37246 6752
rect 37645 6749 37657 6752
rect 37691 6749 37703 6783
rect 37645 6743 37703 6749
rect 34848 6684 34928 6712
rect 34968 6715 35026 6721
rect 34848 6672 34854 6684
rect 34968 6681 34980 6715
rect 35014 6712 35026 6715
rect 36541 6715 36599 6721
rect 36541 6712 36553 6715
rect 35014 6684 36553 6712
rect 35014 6681 35026 6684
rect 34968 6675 35026 6681
rect 36541 6681 36553 6684
rect 36587 6681 36599 6715
rect 36541 6675 36599 6681
rect 31956 6616 32352 6644
rect 33321 6647 33379 6653
rect 33321 6613 33333 6647
rect 33367 6644 33379 6647
rect 33594 6644 33600 6656
rect 33367 6616 33600 6644
rect 33367 6613 33379 6616
rect 33321 6607 33379 6613
rect 33594 6604 33600 6616
rect 33652 6604 33658 6656
rect 35894 6604 35900 6656
rect 35952 6644 35958 6656
rect 36081 6647 36139 6653
rect 36081 6644 36093 6647
rect 35952 6616 36093 6644
rect 35952 6604 35958 6616
rect 36081 6613 36093 6616
rect 36127 6644 36139 6647
rect 36909 6647 36967 6653
rect 36909 6644 36921 6647
rect 36127 6616 36921 6644
rect 36127 6613 36139 6616
rect 36081 6607 36139 6613
rect 36909 6613 36921 6616
rect 36955 6613 36967 6647
rect 36909 6607 36967 6613
rect 37366 6604 37372 6656
rect 37424 6644 37430 6656
rect 37461 6647 37519 6653
rect 37461 6644 37473 6647
rect 37424 6616 37473 6644
rect 37424 6604 37430 6616
rect 37461 6613 37473 6616
rect 37507 6613 37519 6647
rect 37461 6607 37519 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 5626 6440 5632 6452
rect 5539 6412 5632 6440
rect 5626 6400 5632 6412
rect 5684 6440 5690 6452
rect 5810 6440 5816 6452
rect 5684 6412 5816 6440
rect 5684 6400 5690 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 7190 6440 7196 6452
rect 7151 6412 7196 6440
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7834 6440 7840 6452
rect 7760 6412 7840 6440
rect 3694 6372 3700 6384
rect 3160 6344 3700 6372
rect 3160 6313 3188 6344
rect 3694 6332 3700 6344
rect 3752 6332 3758 6384
rect 3878 6332 3884 6384
rect 3936 6332 3942 6384
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4516 6375 4574 6381
rect 4120 6344 4476 6372
rect 4120 6332 4126 6344
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 1872 6100 1900 6267
rect 2516 6236 2544 6267
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3660 6276 3801 6304
rect 3660 6264 3666 6276
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 3896 6304 3924 6332
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 3896 6276 4261 6304
rect 3789 6267 3847 6273
rect 4080 6248 4108 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4448 6304 4476 6344
rect 4516 6341 4528 6375
rect 4562 6372 4574 6375
rect 4706 6372 4712 6384
rect 4562 6344 4712 6372
rect 4562 6341 4574 6344
rect 4516 6335 4574 6341
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 5350 6372 5356 6384
rect 4856 6344 5356 6372
rect 4856 6332 4862 6344
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 7760 6372 7788 6412
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8386 6440 8392 6452
rect 7984 6412 8064 6440
rect 8347 6412 8392 6440
rect 7984 6400 7990 6412
rect 8036 6381 8064 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 11238 6440 11244 6452
rect 9140 6412 11244 6440
rect 6512 6344 7788 6372
rect 8021 6375 8079 6381
rect 6512 6332 6518 6344
rect 8021 6341 8033 6375
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 4448 6276 5672 6304
rect 4249 6267 4307 6273
rect 3878 6236 3884 6248
rect 2516 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 5644 6168 5672 6276
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 5776 6276 6745 6304
rect 5776 6264 5782 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 7006 6304 7012 6316
rect 6967 6276 7012 6304
rect 6733 6267 6791 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 7926 6304 7932 6316
rect 7883 6276 7932 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 8110 6304 8116 6316
rect 8071 6276 8116 6304
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7650 6236 7656 6248
rect 6963 6208 7656 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8220 6236 8248 6267
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8996 6276 9045 6304
rect 8996 6264 9002 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 7800 6208 8248 6236
rect 7800 6196 7806 6208
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9140 6236 9168 6412
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 11974 6440 11980 6452
rect 11747 6412 11980 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 13262 6440 13268 6452
rect 12860 6412 13268 6440
rect 12860 6400 12866 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 15378 6440 15384 6452
rect 15212 6412 15384 6440
rect 9300 6375 9358 6381
rect 9300 6341 9312 6375
rect 9346 6372 9358 6375
rect 10686 6372 10692 6384
rect 9346 6344 9628 6372
rect 9346 6341 9358 6344
rect 9300 6335 9358 6341
rect 9600 6316 9628 6344
rect 10152 6344 10692 6372
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10152 6304 10180 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 11020 6344 13001 6372
rect 11020 6332 11026 6344
rect 12989 6341 13001 6344
rect 13035 6341 13047 6375
rect 12989 6335 13047 6341
rect 13173 6375 13231 6381
rect 13173 6341 13185 6375
rect 13219 6372 13231 6375
rect 13354 6372 13360 6384
rect 13219 6344 13360 6372
rect 13219 6341 13231 6344
rect 13173 6335 13231 6341
rect 13354 6332 13360 6344
rect 13412 6372 13418 6384
rect 13998 6372 14004 6384
rect 13412 6344 14004 6372
rect 13412 6332 13418 6344
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 15102 6372 15108 6384
rect 15063 6344 15108 6372
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 15212 6381 15240 6412
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 15838 6440 15844 6452
rect 15519 6412 15844 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 17037 6443 17095 6449
rect 15988 6412 16033 6440
rect 15988 6400 15994 6412
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17218 6440 17224 6452
rect 17083 6412 17224 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 17310 6400 17316 6452
rect 17368 6400 17374 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 17696 6412 19441 6440
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6341 15255 6375
rect 15562 6372 15568 6384
rect 15197 6335 15255 6341
rect 15304 6344 15568 6372
rect 9732 6276 10180 6304
rect 9732 6264 9738 6276
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 10284 6276 11529 6304
rect 10284 6264 10290 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12618 6304 12624 6316
rect 12483 6276 12624 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 13630 6304 13636 6316
rect 13591 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14550 6304 14556 6316
rect 13955 6276 14556 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 15010 6313 15016 6316
rect 14967 6307 15016 6313
rect 14967 6273 14979 6307
rect 15013 6273 15016 6307
rect 14967 6267 15016 6273
rect 15010 6264 15016 6267
rect 15068 6264 15074 6316
rect 15304 6313 15332 6344
rect 15562 6332 15568 6344
rect 15620 6332 15626 6384
rect 17328 6372 17356 6400
rect 17696 6384 17724 6412
rect 17678 6372 17684 6384
rect 17236 6344 17356 6372
rect 17420 6344 17684 6372
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 15289 6267 15347 6273
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 17236 6313 17264 6344
rect 17222 6307 17280 6313
rect 17222 6273 17234 6307
rect 17268 6273 17280 6307
rect 17222 6267 17280 6273
rect 17313 6307 17371 6313
rect 17313 6273 17325 6307
rect 17359 6304 17371 6307
rect 17420 6304 17448 6344
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 18316 6375 18374 6381
rect 18316 6341 18328 6375
rect 18362 6372 18374 6375
rect 18598 6372 18604 6384
rect 18362 6344 18604 6372
rect 18362 6341 18374 6344
rect 18316 6335 18374 6341
rect 18598 6332 18604 6344
rect 18656 6332 18662 6384
rect 19306 6372 19334 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19978 6440 19984 6452
rect 19939 6412 19984 6440
rect 19429 6403 19487 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20438 6400 20444 6452
rect 20496 6400 20502 6452
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20588 6412 21189 6440
rect 20588 6400 20594 6412
rect 21177 6409 21189 6412
rect 21223 6440 21235 6443
rect 22462 6440 22468 6452
rect 21223 6412 22468 6440
rect 21223 6409 21235 6412
rect 21177 6403 21235 6409
rect 22462 6400 22468 6412
rect 22520 6400 22526 6452
rect 22738 6400 22744 6452
rect 22796 6440 22802 6452
rect 23753 6443 23811 6449
rect 23753 6440 23765 6443
rect 22796 6412 23765 6440
rect 22796 6400 22802 6412
rect 23753 6409 23765 6412
rect 23799 6409 23811 6443
rect 23753 6403 23811 6409
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 24762 6440 24768 6452
rect 24084 6412 24768 6440
rect 24084 6400 24090 6412
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 24854 6400 24860 6452
rect 24912 6440 24918 6452
rect 26237 6443 26295 6449
rect 26237 6440 26249 6443
rect 24912 6412 26249 6440
rect 24912 6400 24918 6412
rect 26237 6409 26249 6412
rect 26283 6409 26295 6443
rect 26237 6403 26295 6409
rect 26878 6400 26884 6452
rect 26936 6440 26942 6452
rect 28353 6443 28411 6449
rect 28353 6440 28365 6443
rect 26936 6412 28365 6440
rect 26936 6400 26942 6412
rect 28353 6409 28365 6412
rect 28399 6409 28411 6443
rect 28353 6403 28411 6409
rect 29641 6443 29699 6449
rect 29641 6409 29653 6443
rect 29687 6440 29699 6443
rect 29730 6440 29736 6452
rect 29687 6412 29736 6440
rect 29687 6409 29699 6412
rect 29641 6403 29699 6409
rect 29730 6400 29736 6412
rect 29788 6400 29794 6452
rect 31846 6400 31852 6452
rect 31904 6440 31910 6452
rect 32769 6443 32827 6449
rect 31904 6412 32720 6440
rect 31904 6400 31910 6412
rect 20456 6372 20484 6400
rect 29270 6372 29276 6384
rect 19306 6344 20484 6372
rect 20548 6344 27972 6372
rect 29231 6344 29276 6372
rect 17586 6304 17592 6316
rect 17359 6276 17448 6304
rect 17547 6276 17592 6304
rect 17359 6273 17371 6276
rect 17313 6267 17371 6273
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 19886 6304 19892 6316
rect 17880 6276 19892 6304
rect 8444 6208 9168 6236
rect 8444 6196 8450 6208
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 12710 6236 12716 6248
rect 11020 6208 12716 6236
rect 11020 6196 11026 6208
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13136 6208 13737 6236
rect 13136 6196 13142 6208
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 17880 6236 17908 6276
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 20036 6276 20177 6304
rect 20036 6264 20042 6276
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20346 6304 20352 6316
rect 20303 6276 20352 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 20548 6313 20576 6344
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20990 6304 20996 6316
rect 20951 6276 20996 6304
rect 20533 6267 20591 6273
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 22094 6304 22100 6316
rect 21324 6276 22100 6304
rect 21324 6264 21330 6276
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 22370 6304 22376 6316
rect 22331 6276 22376 6304
rect 22370 6264 22376 6276
rect 22428 6264 22434 6316
rect 22646 6313 22652 6316
rect 22640 6267 22652 6313
rect 22704 6304 22710 6316
rect 24673 6307 24731 6313
rect 22704 6276 22740 6304
rect 22646 6264 22652 6267
rect 22704 6264 22710 6276
rect 24673 6273 24685 6307
rect 24719 6304 24731 6307
rect 25593 6307 25651 6313
rect 25593 6304 25605 6307
rect 24719 6276 25605 6304
rect 24719 6273 24731 6276
rect 24673 6267 24731 6273
rect 25593 6273 25605 6276
rect 25639 6304 25651 6307
rect 26050 6304 26056 6316
rect 25639 6276 26056 6304
rect 25639 6273 25651 6276
rect 25593 6267 25651 6273
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 26292 6276 26433 6304
rect 26292 6264 26298 6276
rect 26421 6273 26433 6276
rect 26467 6273 26479 6307
rect 26421 6267 26479 6273
rect 26694 6264 26700 6316
rect 26752 6304 26758 6316
rect 27229 6307 27287 6313
rect 27229 6304 27241 6307
rect 26752 6276 27241 6304
rect 26752 6264 26758 6276
rect 27229 6273 27241 6276
rect 27275 6273 27287 6307
rect 27944 6304 27972 6344
rect 29270 6332 29276 6344
rect 29328 6332 29334 6384
rect 29362 6332 29368 6384
rect 29420 6372 29426 6384
rect 29473 6375 29531 6381
rect 29473 6372 29485 6375
rect 29420 6344 29485 6372
rect 29420 6332 29426 6344
rect 29473 6341 29485 6344
rect 29519 6372 29531 6375
rect 31110 6372 31116 6384
rect 29519 6344 31116 6372
rect 29519 6341 29531 6344
rect 29473 6335 29531 6341
rect 27944 6276 28019 6304
rect 27229 6267 27287 6273
rect 18046 6236 18052 6248
rect 13725 6199 13783 6205
rect 15672 6208 17908 6236
rect 18007 6208 18052 6236
rect 8938 6168 8944 6180
rect 2363 6140 4292 6168
rect 5644 6140 8944 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 3418 6100 3424 6112
rect 1872 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3605 6103 3663 6109
rect 3605 6069 3617 6103
rect 3651 6100 3663 6103
rect 3694 6100 3700 6112
rect 3651 6072 3700 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 4264 6100 4292 6140
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11204 6140 12388 6168
rect 11204 6128 11210 6140
rect 5166 6100 5172 6112
rect 4264 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 6454 6100 6460 6112
rect 5500 6072 6460 6100
rect 5500 6060 5506 6072
rect 6454 6060 6460 6072
rect 6512 6060 6518 6112
rect 6730 6100 6736 6112
rect 6691 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 10318 6100 10324 6112
rect 6880 6072 10324 6100
rect 6880 6060 6886 6072
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 10502 6100 10508 6112
rect 10459 6072 10508 6100
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 11848 6072 12265 6100
rect 11848 6060 11854 6072
rect 12253 6069 12265 6072
rect 12299 6069 12311 6103
rect 12360 6100 12388 6140
rect 12618 6128 12624 6180
rect 12676 6168 12682 6180
rect 15672 6168 15700 6208
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 23566 6196 23572 6248
rect 23624 6236 23630 6248
rect 24949 6239 25007 6245
rect 24949 6236 24961 6239
rect 23624 6208 24961 6236
rect 23624 6196 23630 6208
rect 24949 6205 24961 6208
rect 24995 6236 25007 6239
rect 25314 6236 25320 6248
rect 24995 6208 25320 6236
rect 24995 6205 25007 6208
rect 24949 6199 25007 6205
rect 25314 6196 25320 6208
rect 25372 6196 25378 6248
rect 25409 6239 25467 6245
rect 25409 6205 25421 6239
rect 25455 6205 25467 6239
rect 25409 6199 25467 6205
rect 26973 6239 27031 6245
rect 26973 6205 26985 6239
rect 27019 6205 27031 6239
rect 26973 6199 27031 6205
rect 12676 6140 15700 6168
rect 12676 6128 12682 6140
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 15804 6140 18092 6168
rect 15804 6128 15810 6140
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 12360 6072 13645 6100
rect 12253 6063 12311 6069
rect 13633 6069 13645 6072
rect 13679 6069 13691 6103
rect 13633 6063 13691 6069
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14826 6100 14832 6112
rect 14139 6072 14832 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 16666 6100 16672 6112
rect 15068 6072 16672 6100
rect 15068 6060 15074 6072
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17497 6103 17555 6109
rect 17497 6069 17509 6103
rect 17543 6100 17555 6103
rect 17954 6100 17960 6112
rect 17543 6072 17960 6100
rect 17543 6069 17555 6072
rect 17497 6063 17555 6069
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 18064 6100 18092 6140
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 20496 6140 20541 6168
rect 20496 6128 20502 6140
rect 24394 6128 24400 6180
rect 24452 6168 24458 6180
rect 25424 6168 25452 6199
rect 24452 6140 25452 6168
rect 24452 6128 24458 6140
rect 24026 6100 24032 6112
rect 18064 6072 24032 6100
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 24486 6100 24492 6112
rect 24447 6072 24492 6100
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 24857 6103 24915 6109
rect 24857 6069 24869 6103
rect 24903 6100 24915 6103
rect 25130 6100 25136 6112
rect 24903 6072 25136 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 25130 6060 25136 6072
rect 25188 6060 25194 6112
rect 25774 6100 25780 6112
rect 25735 6072 25780 6100
rect 25774 6060 25780 6072
rect 25832 6060 25838 6112
rect 26988 6100 27016 6199
rect 27991 6168 28019 6276
rect 29638 6264 29644 6316
rect 29696 6304 29702 6316
rect 30101 6307 30159 6313
rect 30101 6304 30113 6307
rect 29696 6276 30113 6304
rect 29696 6264 29702 6276
rect 30101 6273 30113 6276
rect 30147 6304 30159 6307
rect 30282 6304 30288 6316
rect 30147 6276 30288 6304
rect 30147 6273 30159 6276
rect 30101 6267 30159 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 30392 6313 30420 6344
rect 31110 6332 31116 6344
rect 31168 6332 31174 6384
rect 32398 6372 32404 6384
rect 32359 6344 32404 6372
rect 32398 6332 32404 6344
rect 32456 6332 32462 6384
rect 32582 6332 32588 6384
rect 32640 6381 32646 6384
rect 32640 6375 32659 6381
rect 32647 6341 32659 6375
rect 32692 6372 32720 6412
rect 32769 6409 32781 6443
rect 32815 6440 32827 6443
rect 32950 6440 32956 6452
rect 32815 6412 32956 6440
rect 32815 6409 32827 6412
rect 32769 6403 32827 6409
rect 32950 6400 32956 6412
rect 33008 6400 33014 6452
rect 33410 6400 33416 6452
rect 33468 6440 33474 6452
rect 34238 6440 34244 6452
rect 33468 6412 34244 6440
rect 33468 6400 33474 6412
rect 34238 6400 34244 6412
rect 34296 6400 34302 6452
rect 36170 6400 36176 6452
rect 36228 6440 36234 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 36228 6412 36553 6440
rect 36228 6400 36234 6412
rect 36541 6409 36553 6412
rect 36587 6409 36599 6443
rect 36541 6403 36599 6409
rect 33226 6372 33232 6384
rect 32692 6344 33232 6372
rect 32640 6335 32659 6341
rect 32640 6332 32646 6335
rect 33226 6332 33232 6344
rect 33284 6332 33290 6384
rect 34146 6332 34152 6384
rect 34204 6372 34210 6384
rect 35428 6375 35486 6381
rect 34204 6344 34928 6372
rect 34204 6332 34210 6344
rect 30377 6307 30435 6313
rect 30377 6273 30389 6307
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 30466 6264 30472 6316
rect 30524 6304 30530 6316
rect 31573 6307 31631 6313
rect 31573 6304 31585 6307
rect 30524 6276 31585 6304
rect 30524 6264 30530 6276
rect 31573 6273 31585 6276
rect 31619 6273 31631 6307
rect 31573 6267 31631 6273
rect 31662 6264 31668 6316
rect 31720 6304 31726 6316
rect 34790 6304 34796 6316
rect 31720 6276 34796 6304
rect 31720 6264 31726 6276
rect 34790 6264 34796 6276
rect 34848 6264 34854 6316
rect 34900 6304 34928 6344
rect 35428 6341 35440 6375
rect 35474 6372 35486 6375
rect 35802 6372 35808 6384
rect 35474 6344 35808 6372
rect 35474 6341 35486 6344
rect 35428 6335 35486 6341
rect 35802 6332 35808 6344
rect 35860 6332 35866 6384
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 34900 6276 37473 6304
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 38105 6307 38163 6313
rect 38105 6273 38117 6307
rect 38151 6273 38163 6307
rect 38105 6267 38163 6273
rect 28074 6196 28080 6248
rect 28132 6236 28138 6248
rect 30834 6236 30840 6248
rect 28132 6208 30840 6236
rect 28132 6196 28138 6208
rect 30834 6196 30840 6208
rect 30892 6196 30898 6248
rect 31202 6196 31208 6248
rect 31260 6236 31266 6248
rect 33321 6239 33379 6245
rect 31260 6208 33272 6236
rect 31260 6196 31266 6208
rect 32490 6168 32496 6180
rect 27991 6140 32496 6168
rect 32490 6128 32496 6140
rect 32548 6128 32554 6180
rect 33244 6168 33272 6208
rect 33321 6205 33333 6239
rect 33367 6236 33379 6239
rect 33410 6236 33416 6248
rect 33367 6208 33416 6236
rect 33367 6205 33379 6208
rect 33321 6199 33379 6205
rect 33410 6196 33416 6208
rect 33468 6196 33474 6248
rect 33597 6239 33655 6245
rect 33597 6205 33609 6239
rect 33643 6205 33655 6239
rect 33597 6199 33655 6205
rect 33612 6168 33640 6199
rect 34698 6196 34704 6248
rect 34756 6236 34762 6248
rect 35161 6239 35219 6245
rect 35161 6236 35173 6239
rect 34756 6208 35173 6236
rect 34756 6196 34762 6208
rect 35161 6205 35173 6208
rect 35207 6205 35219 6239
rect 35161 6199 35219 6205
rect 36814 6196 36820 6248
rect 36872 6236 36878 6248
rect 38120 6236 38148 6267
rect 36872 6208 38148 6236
rect 36872 6196 36878 6208
rect 34330 6168 34336 6180
rect 33244 6140 34336 6168
rect 34330 6128 34336 6140
rect 34388 6128 34394 6180
rect 28166 6100 28172 6112
rect 26988 6072 28172 6100
rect 28166 6060 28172 6072
rect 28224 6060 28230 6112
rect 28258 6060 28264 6112
rect 28316 6100 28322 6112
rect 28718 6100 28724 6112
rect 28316 6072 28724 6100
rect 28316 6060 28322 6072
rect 28718 6060 28724 6072
rect 28776 6060 28782 6112
rect 29454 6100 29460 6112
rect 29415 6072 29460 6100
rect 29454 6060 29460 6072
rect 29512 6060 29518 6112
rect 29730 6060 29736 6112
rect 29788 6100 29794 6112
rect 30098 6100 30104 6112
rect 29788 6072 30104 6100
rect 29788 6060 29794 6072
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 31018 6060 31024 6112
rect 31076 6100 31082 6112
rect 31389 6103 31447 6109
rect 31389 6100 31401 6103
rect 31076 6072 31401 6100
rect 31076 6060 31082 6072
rect 31389 6069 31401 6072
rect 31435 6069 31447 6103
rect 31389 6063 31447 6069
rect 32585 6103 32643 6109
rect 32585 6069 32597 6103
rect 32631 6100 32643 6103
rect 33778 6100 33784 6112
rect 32631 6072 33784 6100
rect 32631 6069 32643 6072
rect 32585 6063 32643 6069
rect 33778 6060 33784 6072
rect 33836 6100 33842 6112
rect 34422 6100 34428 6112
rect 33836 6072 34428 6100
rect 33836 6060 33842 6072
rect 34422 6060 34428 6072
rect 34480 6060 34486 6112
rect 36354 6060 36360 6112
rect 36412 6100 36418 6112
rect 37277 6103 37335 6109
rect 37277 6100 37289 6103
rect 36412 6072 37289 6100
rect 36412 6060 36418 6072
rect 37277 6069 37289 6072
rect 37323 6069 37335 6103
rect 37277 6063 37335 6069
rect 37458 6060 37464 6112
rect 37516 6100 37522 6112
rect 37921 6103 37979 6109
rect 37921 6100 37933 6103
rect 37516 6072 37933 6100
rect 37516 6060 37522 6072
rect 37921 6069 37933 6072
rect 37967 6069 37979 6103
rect 37921 6063 37979 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 5534 5896 5540 5908
rect 1811 5868 5396 5896
rect 5495 5868 5540 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 3694 5828 3700 5840
rect 2455 5800 3700 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 3694 5788 3700 5800
rect 3752 5788 3758 5840
rect 5368 5828 5396 5868
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 10962 5896 10968 5908
rect 5644 5868 10968 5896
rect 5644 5828 5672 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11974 5896 11980 5908
rect 11388 5868 11980 5896
rect 11388 5856 11394 5868
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12342 5896 12348 5908
rect 12303 5868 12348 5896
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 15010 5896 15016 5908
rect 14700 5868 15016 5896
rect 14700 5856 14706 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15194 5896 15200 5908
rect 15151 5868 15200 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 18601 5899 18659 5905
rect 18601 5896 18613 5899
rect 16172 5868 18613 5896
rect 16172 5856 16178 5868
rect 18601 5865 18613 5868
rect 18647 5865 18659 5899
rect 18601 5859 18659 5865
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20404 5868 21005 5896
rect 20404 5856 20410 5868
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 23382 5896 23388 5908
rect 21039 5868 23388 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23532 5868 23577 5896
rect 23532 5856 23538 5868
rect 25314 5856 25320 5908
rect 25372 5896 25378 5908
rect 25777 5899 25835 5905
rect 25777 5896 25789 5899
rect 25372 5868 25789 5896
rect 25372 5856 25378 5868
rect 25777 5865 25789 5868
rect 25823 5865 25835 5899
rect 25777 5859 25835 5865
rect 26050 5856 26056 5908
rect 26108 5896 26114 5908
rect 27617 5899 27675 5905
rect 26108 5868 27568 5896
rect 26108 5856 26114 5868
rect 5368 5800 5672 5828
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8662 5828 8668 5840
rect 8435 5800 8668 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 13541 5831 13599 5837
rect 8996 5800 10548 5828
rect 8996 5788 9002 5800
rect 3142 5760 3148 5772
rect 2608 5732 3148 5760
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2498 5692 2504 5704
rect 1995 5664 2504 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2608 5701 2636 5732
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 4120 5732 4169 5760
rect 4120 5720 4126 5732
rect 4157 5729 4169 5732
rect 4203 5729 4215 5763
rect 4157 5723 4215 5729
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 5868 5732 10425 5760
rect 5868 5720 5874 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 3283 5664 6377 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 9122 5692 9128 5704
rect 7515 5664 9128 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 9232 5664 9321 5692
rect 4402 5627 4460 5633
rect 4402 5624 4414 5627
rect 3068 5596 4414 5624
rect 3068 5565 3096 5596
rect 4402 5593 4414 5596
rect 4448 5593 4460 5627
rect 4402 5587 4460 5593
rect 5258 5584 5264 5636
rect 5316 5624 5322 5636
rect 5997 5627 6055 5633
rect 5997 5624 6009 5627
rect 5316 5596 6009 5624
rect 5316 5584 5322 5596
rect 5997 5593 6009 5596
rect 6043 5593 6055 5627
rect 5997 5587 6055 5593
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 6181 5627 6239 5633
rect 6181 5624 6193 5627
rect 6144 5596 6193 5624
rect 6144 5584 6150 5596
rect 6181 5593 6193 5596
rect 6227 5593 6239 5627
rect 6181 5587 6239 5593
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 7248 5596 8156 5624
rect 7248 5584 7254 5596
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5525 3111 5559
rect 3053 5519 3111 5525
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 5074 5556 5080 5568
rect 3936 5528 5080 5556
rect 3936 5516 3942 5528
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 6972 5528 7573 5556
rect 6972 5516 6978 5528
rect 7561 5525 7573 5528
rect 7607 5525 7619 5559
rect 8128 5556 8156 5596
rect 8202 5584 8208 5636
rect 8260 5624 8266 5636
rect 8260 5596 8305 5624
rect 8260 5584 8266 5596
rect 9232 5556 9260 5664
rect 9309 5661 9321 5664
rect 9355 5692 9367 5695
rect 10226 5692 10232 5704
rect 9355 5664 10232 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10137 5627 10195 5633
rect 10137 5593 10149 5627
rect 10183 5593 10195 5627
rect 10137 5587 10195 5593
rect 9490 5556 9496 5568
rect 8128 5528 9260 5556
rect 9451 5528 9496 5556
rect 7561 5519 7619 5525
rect 9490 5516 9496 5528
rect 9548 5556 9554 5568
rect 10042 5556 10048 5568
rect 9548 5528 10048 5556
rect 9548 5516 9554 5528
rect 10042 5516 10048 5528
rect 10100 5556 10106 5568
rect 10152 5556 10180 5587
rect 10100 5528 10180 5556
rect 10428 5556 10456 5723
rect 10520 5624 10548 5800
rect 13541 5797 13553 5831
rect 13587 5828 13599 5831
rect 14182 5828 14188 5840
rect 13587 5800 14188 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 12526 5760 12532 5772
rect 11983 5732 12532 5760
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11983 5692 12011 5732
rect 12526 5720 12532 5732
rect 12584 5760 12590 5772
rect 13556 5760 13584 5791
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 14918 5788 14924 5840
rect 14976 5828 14982 5840
rect 14976 5800 15332 5828
rect 14976 5788 14982 5800
rect 15102 5760 15108 5772
rect 12584 5732 13584 5760
rect 15063 5732 15108 5760
rect 12584 5720 12590 5732
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15304 5760 15332 5800
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 16942 5828 16948 5840
rect 15804 5800 16948 5828
rect 15804 5788 15810 5800
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17681 5831 17739 5837
rect 17681 5797 17693 5831
rect 17727 5828 17739 5831
rect 22465 5831 22523 5837
rect 22465 5828 22477 5831
rect 17727 5800 17908 5828
rect 17727 5797 17739 5800
rect 17681 5791 17739 5797
rect 16114 5760 16120 5772
rect 15304 5732 16120 5760
rect 13354 5692 13360 5704
rect 11011 5664 12011 5692
rect 13315 5664 13360 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 15304 5701 15332 5732
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16850 5760 16856 5772
rect 16224 5732 16856 5760
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 15289 5695 15347 5701
rect 14415 5664 15240 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 11210 5627 11268 5633
rect 11210 5624 11222 5627
rect 10520 5596 11222 5624
rect 11210 5593 11222 5596
rect 11256 5593 11268 5627
rect 14182 5624 14188 5636
rect 11210 5587 11268 5593
rect 11348 5596 14188 5624
rect 11348 5556 11376 5596
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 14550 5624 14556 5636
rect 14511 5596 14556 5624
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 14918 5584 14924 5636
rect 14976 5624 14982 5636
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 14976 5596 15025 5624
rect 14976 5584 14982 5596
rect 15013 5593 15025 5596
rect 15059 5593 15071 5627
rect 15212 5624 15240 5664
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 16224 5701 16252 5732
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 17276 5732 17448 5760
rect 17276 5720 17282 5732
rect 16209 5695 16267 5701
rect 16209 5692 16221 5695
rect 15436 5664 16221 5692
rect 15436 5652 15442 5664
rect 16209 5661 16221 5664
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 16574 5692 16580 5704
rect 16531 5664 16580 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 17420 5701 17448 5732
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17880 5760 17908 5800
rect 22066 5800 22477 5828
rect 17954 5760 17960 5772
rect 17644 5732 17816 5760
rect 17880 5732 17960 5760
rect 17644 5720 17650 5732
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17678 5692 17684 5704
rect 17543 5664 17684 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 17788 5701 17816 5732
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 19613 5763 19671 5769
rect 19613 5760 19625 5763
rect 18104 5732 19625 5760
rect 18104 5720 18110 5732
rect 19613 5729 19625 5732
rect 19659 5729 19671 5763
rect 22066 5760 22094 5800
rect 22465 5797 22477 5800
rect 22511 5828 22523 5831
rect 22738 5828 22744 5840
rect 22511 5800 22744 5828
rect 22511 5797 22523 5800
rect 22465 5791 22523 5797
rect 22738 5788 22744 5800
rect 22796 5788 22802 5840
rect 27540 5828 27568 5868
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27798 5896 27804 5908
rect 27663 5868 27804 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 27798 5856 27804 5868
rect 27856 5856 27862 5908
rect 29454 5856 29460 5908
rect 29512 5896 29518 5908
rect 29917 5899 29975 5905
rect 29917 5896 29929 5899
rect 29512 5868 29929 5896
rect 29512 5856 29518 5868
rect 29917 5865 29929 5868
rect 29963 5896 29975 5899
rect 31202 5896 31208 5908
rect 29963 5868 31208 5896
rect 29963 5865 29975 5868
rect 29917 5859 29975 5865
rect 31202 5856 31208 5868
rect 31260 5856 31266 5908
rect 31754 5856 31760 5908
rect 31812 5896 31818 5908
rect 32953 5899 33011 5905
rect 32953 5896 32965 5899
rect 31812 5868 32965 5896
rect 31812 5856 31818 5868
rect 32953 5865 32965 5868
rect 32999 5865 33011 5899
rect 33778 5896 33784 5908
rect 33739 5868 33784 5896
rect 32953 5859 33011 5865
rect 33778 5856 33784 5868
rect 33836 5856 33842 5908
rect 33870 5856 33876 5908
rect 33928 5896 33934 5908
rect 33965 5899 34023 5905
rect 33965 5896 33977 5899
rect 33928 5868 33977 5896
rect 33928 5856 33934 5868
rect 33965 5865 33977 5868
rect 34011 5865 34023 5899
rect 33965 5859 34023 5865
rect 34422 5856 34428 5908
rect 34480 5896 34486 5908
rect 34606 5896 34612 5908
rect 34480 5868 34612 5896
rect 34480 5856 34486 5868
rect 34606 5856 34612 5868
rect 34664 5896 34670 5908
rect 35161 5899 35219 5905
rect 35161 5896 35173 5899
rect 34664 5868 35173 5896
rect 34664 5856 34670 5868
rect 35161 5865 35173 5868
rect 35207 5865 35219 5899
rect 35161 5859 35219 5865
rect 35345 5899 35403 5905
rect 35345 5865 35357 5899
rect 35391 5896 35403 5899
rect 36446 5896 36452 5908
rect 35391 5868 36452 5896
rect 35391 5865 35403 5868
rect 35345 5859 35403 5865
rect 36446 5856 36452 5868
rect 36504 5856 36510 5908
rect 29362 5828 29368 5840
rect 27540 5800 29368 5828
rect 29362 5788 29368 5800
rect 29420 5788 29426 5840
rect 30006 5788 30012 5840
rect 30064 5828 30070 5840
rect 30101 5831 30159 5837
rect 30101 5828 30113 5831
rect 30064 5800 30113 5828
rect 30064 5788 30070 5800
rect 30101 5797 30113 5800
rect 30147 5797 30159 5831
rect 30374 5828 30380 5840
rect 30101 5791 30159 5797
rect 30208 5800 30380 5828
rect 23566 5760 23572 5772
rect 19613 5723 19671 5729
rect 20640 5732 22094 5760
rect 22848 5732 23572 5760
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 18414 5692 18420 5704
rect 18375 5664 18420 5692
rect 17773 5655 17831 5661
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19869 5695 19927 5701
rect 19869 5692 19881 5695
rect 19392 5664 19881 5692
rect 19392 5652 19398 5664
rect 19869 5661 19881 5664
rect 19915 5661 19927 5695
rect 19869 5655 19927 5661
rect 15930 5624 15936 5636
rect 15212 5596 15936 5624
rect 15013 5587 15071 5593
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 16025 5627 16083 5633
rect 16025 5624 16037 5627
rect 15988 5596 16037 5624
rect 15988 5584 15994 5596
rect 16025 5593 16037 5596
rect 16071 5593 16083 5627
rect 16025 5587 16083 5593
rect 17221 5627 17279 5633
rect 17221 5593 17233 5627
rect 17267 5624 17279 5627
rect 18233 5627 18291 5633
rect 18233 5624 18245 5627
rect 17267 5596 18245 5624
rect 17267 5593 17279 5596
rect 17221 5587 17279 5593
rect 18233 5593 18245 5596
rect 18279 5593 18291 5627
rect 18233 5587 18291 5593
rect 10428 5528 11376 5556
rect 10100 5516 10106 5528
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 13688 5528 15485 5556
rect 13688 5516 13694 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 15473 5519 15531 5525
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 17034 5556 17040 5568
rect 16439 5528 17040 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 17034 5516 17040 5528
rect 17092 5556 17098 5568
rect 20640 5556 20668 5732
rect 22002 5692 22008 5704
rect 21963 5664 22008 5692
rect 22002 5652 22008 5664
rect 22060 5692 22066 5704
rect 22848 5692 22876 5732
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 27430 5720 27436 5772
rect 27488 5760 27494 5772
rect 30208 5760 30236 5800
rect 30374 5788 30380 5800
rect 30432 5788 30438 5840
rect 33137 5831 33195 5837
rect 33137 5797 33149 5831
rect 33183 5828 33195 5831
rect 33183 5800 37320 5828
rect 33183 5797 33195 5800
rect 33137 5791 33195 5797
rect 27488 5732 30236 5760
rect 27488 5720 27494 5732
rect 30282 5720 30288 5772
rect 30340 5760 30346 5772
rect 31481 5763 31539 5769
rect 31481 5760 31493 5763
rect 30340 5732 31493 5760
rect 30340 5720 30346 5732
rect 31481 5729 31493 5732
rect 31527 5729 31539 5763
rect 31481 5723 31539 5729
rect 31757 5763 31815 5769
rect 31757 5729 31769 5763
rect 31803 5760 31815 5763
rect 32582 5760 32588 5772
rect 31803 5732 32588 5760
rect 31803 5729 31815 5732
rect 31757 5723 31815 5729
rect 32582 5720 32588 5732
rect 32640 5720 32646 5772
rect 22060 5664 22876 5692
rect 22060 5652 22066 5664
rect 22922 5652 22928 5704
rect 22980 5692 22986 5704
rect 23293 5695 23351 5701
rect 23293 5692 23305 5695
rect 22980 5664 23305 5692
rect 22980 5652 22986 5664
rect 23293 5661 23305 5664
rect 23339 5692 23351 5695
rect 23382 5692 23388 5704
rect 23339 5664 23388 5692
rect 23339 5661 23351 5664
rect 23293 5655 23351 5661
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 24302 5652 24308 5704
rect 24360 5692 24366 5704
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 24360 5664 24409 5692
rect 24360 5652 24366 5664
rect 24397 5661 24409 5664
rect 24443 5692 24455 5695
rect 26237 5695 26295 5701
rect 26237 5692 26249 5695
rect 24443 5664 26249 5692
rect 24443 5661 24455 5664
rect 24397 5655 24455 5661
rect 26237 5661 26249 5664
rect 26283 5692 26295 5695
rect 27522 5692 27528 5704
rect 26283 5664 27528 5692
rect 26283 5661 26295 5664
rect 26237 5655 26295 5661
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 28353 5695 28411 5701
rect 28353 5692 28365 5695
rect 27764 5664 28365 5692
rect 27764 5652 27770 5664
rect 28353 5661 28365 5664
rect 28399 5692 28411 5695
rect 28810 5692 28816 5704
rect 28399 5664 28816 5692
rect 28399 5661 28411 5664
rect 28353 5655 28411 5661
rect 28810 5652 28816 5664
rect 28868 5652 28874 5704
rect 28994 5692 29000 5704
rect 28955 5664 29000 5692
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 29362 5652 29368 5704
rect 29420 5692 29426 5704
rect 30742 5692 30748 5704
rect 29420 5664 29960 5692
rect 30703 5664 30748 5692
rect 29420 5652 29426 5664
rect 24486 5584 24492 5636
rect 24544 5624 24550 5636
rect 24642 5627 24700 5633
rect 24642 5624 24654 5627
rect 24544 5596 24654 5624
rect 24544 5584 24550 5596
rect 24642 5593 24654 5596
rect 24688 5593 24700 5627
rect 24642 5587 24700 5593
rect 26504 5627 26562 5633
rect 26504 5593 26516 5627
rect 26550 5624 26562 5627
rect 26878 5624 26884 5636
rect 26550 5596 26884 5624
rect 26550 5593 26562 5596
rect 26504 5587 26562 5593
rect 26878 5584 26884 5596
rect 26936 5584 26942 5636
rect 26970 5584 26976 5636
rect 27028 5624 27034 5636
rect 29733 5627 29791 5633
rect 27028 5596 28856 5624
rect 27028 5584 27034 5596
rect 17092 5528 20668 5556
rect 17092 5516 17098 5528
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 22005 5559 22063 5565
rect 22005 5556 22017 5559
rect 21784 5528 22017 5556
rect 21784 5516 21790 5528
rect 22005 5525 22017 5528
rect 22051 5525 22063 5559
rect 22005 5519 22063 5525
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23290 5556 23296 5568
rect 22796 5528 23296 5556
rect 22796 5516 22802 5528
rect 23290 5516 23296 5528
rect 23348 5516 23354 5568
rect 23658 5516 23664 5568
rect 23716 5556 23722 5568
rect 23845 5559 23903 5565
rect 23845 5556 23857 5559
rect 23716 5528 23857 5556
rect 23716 5516 23722 5528
rect 23845 5525 23857 5528
rect 23891 5525 23903 5559
rect 23845 5519 23903 5525
rect 28169 5559 28227 5565
rect 28169 5525 28181 5559
rect 28215 5556 28227 5559
rect 28718 5556 28724 5568
rect 28215 5528 28724 5556
rect 28215 5525 28227 5528
rect 28169 5519 28227 5525
rect 28718 5516 28724 5528
rect 28776 5516 28782 5568
rect 28828 5565 28856 5596
rect 29733 5593 29745 5627
rect 29779 5624 29791 5627
rect 29822 5624 29828 5636
rect 29779 5596 29828 5624
rect 29779 5593 29791 5596
rect 29733 5587 29791 5593
rect 29822 5584 29828 5596
rect 29880 5584 29886 5636
rect 29932 5633 29960 5664
rect 30742 5652 30748 5664
rect 30800 5652 30806 5704
rect 29932 5627 29991 5633
rect 29932 5596 29945 5627
rect 29933 5593 29945 5596
rect 29979 5593 29991 5627
rect 31294 5624 31300 5636
rect 29933 5587 29991 5593
rect 30024 5596 31300 5624
rect 28813 5559 28871 5565
rect 28813 5525 28825 5559
rect 28859 5525 28871 5559
rect 28813 5519 28871 5525
rect 28902 5516 28908 5568
rect 28960 5556 28966 5568
rect 30024 5556 30052 5596
rect 31294 5584 31300 5596
rect 31352 5584 31358 5636
rect 28960 5528 30052 5556
rect 28960 5516 28966 5528
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 30561 5559 30619 5565
rect 30561 5556 30573 5559
rect 30432 5528 30573 5556
rect 30432 5516 30438 5528
rect 30561 5525 30573 5528
rect 30607 5525 30619 5559
rect 32600 5556 32628 5720
rect 32876 5664 33180 5692
rect 32769 5627 32827 5633
rect 32769 5593 32781 5627
rect 32815 5624 32827 5627
rect 32876 5624 32904 5664
rect 32815 5596 32904 5624
rect 32815 5593 32827 5596
rect 32769 5587 32827 5593
rect 32950 5584 32956 5636
rect 33008 5633 33014 5636
rect 33008 5627 33027 5633
rect 33015 5593 33027 5627
rect 33152 5624 33180 5664
rect 33226 5652 33232 5704
rect 33284 5692 33290 5704
rect 35820 5701 36008 5708
rect 35820 5695 36047 5701
rect 35820 5692 36001 5695
rect 33284 5680 36001 5692
rect 33284 5664 35848 5680
rect 35980 5664 36001 5680
rect 33284 5652 33290 5664
rect 35989 5661 36001 5664
rect 36035 5661 36047 5695
rect 35989 5655 36047 5661
rect 36078 5652 36084 5704
rect 36136 5692 36142 5704
rect 37292 5701 37320 5800
rect 36633 5695 36691 5701
rect 36633 5692 36645 5695
rect 36136 5664 36645 5692
rect 36136 5652 36142 5664
rect 36633 5661 36645 5664
rect 36679 5661 36691 5695
rect 36633 5655 36691 5661
rect 37277 5695 37335 5701
rect 37277 5661 37289 5695
rect 37323 5661 37335 5695
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37277 5655 37335 5661
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 33594 5624 33600 5636
rect 33152 5596 33600 5624
rect 33008 5587 33027 5593
rect 33008 5584 33014 5587
rect 33594 5584 33600 5596
rect 33652 5584 33658 5636
rect 34977 5627 35035 5633
rect 34977 5593 34989 5627
rect 35023 5624 35035 5627
rect 36538 5624 36544 5636
rect 35023 5596 36544 5624
rect 35023 5593 35035 5596
rect 34977 5587 35035 5593
rect 36538 5584 36544 5596
rect 36596 5584 36602 5636
rect 33797 5559 33855 5565
rect 33797 5556 33809 5559
rect 32600 5528 33809 5556
rect 30561 5519 30619 5525
rect 33797 5525 33809 5528
rect 33843 5556 33855 5559
rect 34790 5556 34796 5568
rect 33843 5528 34796 5556
rect 33843 5525 33855 5528
rect 33797 5519 33855 5525
rect 34790 5516 34796 5528
rect 34848 5556 34854 5568
rect 35177 5559 35235 5565
rect 35177 5556 35189 5559
rect 34848 5528 35189 5556
rect 34848 5516 34854 5528
rect 35177 5525 35189 5528
rect 35223 5525 35235 5559
rect 35177 5519 35235 5525
rect 35526 5516 35532 5568
rect 35584 5556 35590 5568
rect 35805 5559 35863 5565
rect 35805 5556 35817 5559
rect 35584 5528 35817 5556
rect 35584 5516 35590 5528
rect 35805 5525 35817 5528
rect 35851 5525 35863 5559
rect 35805 5519 35863 5525
rect 35986 5516 35992 5568
rect 36044 5556 36050 5568
rect 36449 5559 36507 5565
rect 36449 5556 36461 5559
rect 36044 5528 36461 5556
rect 36044 5516 36050 5528
rect 36449 5525 36461 5528
rect 36495 5525 36507 5559
rect 37090 5556 37096 5568
rect 37051 5528 37096 5556
rect 36449 5519 36507 5525
rect 37090 5516 37096 5528
rect 37148 5516 37154 5568
rect 38013 5559 38071 5565
rect 38013 5525 38025 5559
rect 38059 5556 38071 5559
rect 39390 5556 39396 5568
rect 38059 5528 39396 5556
rect 38059 5525 38071 5528
rect 38013 5519 38071 5525
rect 39390 5516 39396 5528
rect 39448 5516 39454 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 2363 5324 4844 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 4062 5284 4068 5296
rect 2976 5256 4068 5284
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2498 5216 2504 5228
rect 2459 5188 2504 5216
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2976 5225 3004 5256
rect 4062 5244 4068 5256
rect 4120 5284 4126 5296
rect 4614 5284 4620 5296
rect 4120 5256 4620 5284
rect 4120 5244 4126 5256
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 4816 5284 4844 5324
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 4948 5324 5181 5352
rect 4948 5312 4954 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 5169 5315 5227 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8168 5324 8309 5352
rect 8168 5312 8174 5324
rect 8297 5321 8309 5324
rect 8343 5352 8355 5355
rect 9030 5352 9036 5364
rect 8343 5324 9036 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9677 5355 9735 5361
rect 9677 5321 9689 5355
rect 9723 5352 9735 5355
rect 10134 5352 10140 5364
rect 9723 5324 10140 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 10376 5324 11897 5352
rect 10376 5312 10382 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 13538 5352 13544 5364
rect 12032 5324 13544 5352
rect 12032 5312 12038 5324
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 14090 5352 14096 5364
rect 13955 5324 14096 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 19426 5352 19432 5364
rect 15764 5324 19432 5352
rect 7184 5287 7242 5293
rect 4816 5256 7144 5284
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3217 5219 3275 5225
rect 3217 5216 3229 5219
rect 3108 5188 3229 5216
rect 3108 5176 3114 5188
rect 3217 5185 3229 5188
rect 3263 5185 3275 5219
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 3217 5179 3275 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 5810 5216 5816 5228
rect 5771 5188 5816 5216
rect 4985 5179 5043 5185
rect 5000 5148 5028 5179
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6914 5216 6920 5228
rect 6512 5188 6920 5216
rect 6512 5176 6518 5188
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7116 5216 7144 5256
rect 7184 5253 7196 5287
rect 7230 5284 7242 5287
rect 7374 5284 7380 5296
rect 7230 5256 7380 5284
rect 7230 5253 7242 5256
rect 7184 5247 7242 5253
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 8662 5244 8668 5296
rect 8720 5284 8726 5296
rect 9493 5287 9551 5293
rect 9493 5284 9505 5287
rect 8720 5256 9505 5284
rect 8720 5244 8726 5256
rect 9493 5253 9505 5256
rect 9539 5253 9551 5287
rect 9493 5247 9551 5253
rect 7466 5216 7472 5228
rect 7116 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 9306 5216 9312 5228
rect 9267 5188 9312 5216
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9508 5216 9536 5247
rect 9766 5244 9772 5296
rect 9824 5284 9830 5296
rect 10870 5284 10876 5296
rect 9824 5256 10876 5284
rect 9824 5244 9830 5256
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 12774 5287 12832 5293
rect 12774 5284 12786 5287
rect 11072 5256 12786 5284
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9508 5188 10425 5216
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 4264 5120 5028 5148
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4264 5012 4292 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10100 5120 10149 5148
rect 10100 5108 10106 5120
rect 10137 5117 10149 5120
rect 10183 5148 10195 5151
rect 10962 5148 10968 5160
rect 10183 5120 10968 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 4706 5080 4712 5092
rect 4387 5052 4712 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 4706 5040 4712 5052
rect 4764 5080 4770 5092
rect 5718 5080 5724 5092
rect 4764 5052 5724 5080
rect 4764 5040 4770 5052
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 11072 5080 11100 5256
rect 12774 5253 12786 5256
rect 12820 5253 12832 5287
rect 15378 5284 15384 5296
rect 12774 5247 12832 5253
rect 14568 5256 15384 5284
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11422 5216 11428 5228
rect 11204 5188 11428 5216
rect 11204 5176 11210 5188
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11606 5216 11612 5228
rect 11563 5188 11612 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 8352 5052 11100 5080
rect 11716 5080 11744 5179
rect 12526 5176 12532 5228
rect 12584 5225 12590 5228
rect 12584 5216 12594 5225
rect 12584 5188 12629 5216
rect 12584 5179 12594 5188
rect 12584 5176 12590 5179
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 14568 5216 14596 5256
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 15102 5216 15108 5228
rect 13136 5188 14596 5216
rect 15063 5188 15108 5216
rect 13136 5176 13142 5188
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15473 5219 15531 5225
rect 15252 5188 15297 5216
rect 15252 5176 15258 5188
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 15764 5216 15792 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 22554 5312 22560 5364
rect 22612 5352 22618 5364
rect 22833 5355 22891 5361
rect 22833 5352 22845 5355
rect 22612 5324 22845 5352
rect 22612 5312 22618 5324
rect 22833 5321 22845 5324
rect 22879 5321 22891 5355
rect 22833 5315 22891 5321
rect 24121 5355 24179 5361
rect 24121 5321 24133 5355
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 24412 5324 27844 5352
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 15948 5256 17049 5284
rect 15948 5228 15976 5256
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 24136 5284 24164 5315
rect 17037 5247 17095 5253
rect 19720 5256 24164 5284
rect 15930 5216 15936 5228
rect 15519 5188 15792 5216
rect 15891 5188 15936 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16482 5216 16488 5228
rect 16163 5188 16488 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 18966 5216 18972 5228
rect 18927 5188 18972 5216
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19720 5225 19748 5256
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5185 19763 5219
rect 20714 5216 20720 5228
rect 20675 5188 20720 5216
rect 19705 5179 19763 5185
rect 20714 5176 20720 5188
rect 20772 5216 20778 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 20772 5188 21833 5216
rect 20772 5176 20778 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22005 5219 22063 5225
rect 22005 5185 22017 5219
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22278 5216 22284 5228
rect 22235 5188 22284 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 15286 5148 15292 5160
rect 13964 5120 15292 5148
rect 13964 5108 13970 5120
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15436 5120 16037 5148
rect 15436 5108 15442 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 17681 5151 17739 5157
rect 17681 5148 17693 5151
rect 16025 5111 16083 5117
rect 17144 5120 17693 5148
rect 12526 5080 12532 5092
rect 11716 5052 12532 5080
rect 8352 5040 8358 5052
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 4120 4984 5641 5012
rect 4120 4972 4126 4984
rect 5629 4981 5641 4984
rect 5675 5012 5687 5015
rect 6086 5012 6092 5024
rect 5675 4984 6092 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 11716 5012 11744 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 6420 4984 11744 5012
rect 14921 5015 14979 5021
rect 6420 4972 6426 4984
rect 14921 4981 14933 5015
rect 14967 5012 14979 5015
rect 15286 5012 15292 5024
rect 14967 4984 15292 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 15381 5015 15439 5021
rect 15381 4981 15393 5015
rect 15427 5012 15439 5015
rect 15470 5012 15476 5024
rect 15427 4984 15476 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 15470 4972 15476 4984
rect 15528 5012 15534 5024
rect 17144 5021 17172 5120
rect 17681 5117 17693 5120
rect 17727 5117 17739 5151
rect 17954 5148 17960 5160
rect 17867 5120 17960 5148
rect 17681 5111 17739 5117
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 22020 5148 22048 5179
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 22738 5216 22744 5228
rect 22695 5188 22744 5216
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 22925 5220 22983 5225
rect 22925 5219 23000 5220
rect 22925 5185 22937 5219
rect 22971 5185 23000 5219
rect 22925 5179 23000 5185
rect 22972 5148 23000 5179
rect 23290 5176 23296 5228
rect 23348 5216 23354 5228
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 23348 5188 23397 5216
rect 23348 5176 23354 5188
rect 23385 5185 23397 5188
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 23569 5219 23627 5225
rect 23569 5185 23581 5219
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23584 5148 23612 5179
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 24302 5216 24308 5228
rect 23716 5188 23761 5216
rect 24263 5188 24308 5216
rect 23716 5176 23722 5188
rect 24302 5176 24308 5188
rect 24360 5176 24366 5228
rect 20864 5120 22048 5148
rect 22112 5120 23612 5148
rect 20864 5108 20870 5120
rect 17972 5080 18000 5108
rect 20438 5080 20444 5092
rect 17972 5052 20444 5080
rect 20438 5040 20444 5052
rect 20496 5080 20502 5092
rect 22112 5080 22140 5120
rect 24026 5108 24032 5160
rect 24084 5148 24090 5160
rect 24412 5148 24440 5324
rect 25314 5244 25320 5296
rect 25372 5284 25378 5296
rect 27706 5284 27712 5296
rect 25372 5256 27712 5284
rect 25372 5244 25378 5256
rect 27706 5244 27712 5256
rect 27764 5244 27770 5296
rect 24946 5216 24952 5228
rect 24859 5188 24952 5216
rect 24946 5176 24952 5188
rect 25004 5216 25010 5228
rect 25590 5216 25596 5228
rect 25004 5188 25452 5216
rect 25551 5188 25596 5216
rect 25004 5176 25010 5188
rect 24084 5120 24440 5148
rect 25424 5148 25452 5188
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 25682 5176 25688 5228
rect 25740 5216 25746 5228
rect 26237 5219 26295 5225
rect 26237 5216 26249 5219
rect 25740 5188 26249 5216
rect 25740 5176 25746 5188
rect 26237 5185 26249 5188
rect 26283 5185 26295 5219
rect 26237 5179 26295 5185
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27816 5216 27844 5324
rect 28902 5312 28908 5364
rect 28960 5352 28966 5364
rect 29381 5355 29439 5361
rect 29381 5352 29393 5355
rect 28960 5324 29393 5352
rect 28960 5312 28966 5324
rect 29381 5321 29393 5324
rect 29427 5352 29439 5355
rect 29549 5355 29607 5361
rect 29427 5324 29500 5352
rect 29427 5321 29439 5324
rect 29381 5315 29439 5321
rect 28261 5287 28319 5293
rect 28261 5253 28273 5287
rect 28307 5284 28319 5287
rect 28534 5284 28540 5296
rect 28307 5256 28540 5284
rect 28307 5253 28319 5256
rect 28261 5247 28319 5253
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 29181 5287 29239 5293
rect 29181 5253 29193 5287
rect 29227 5284 29239 5287
rect 29270 5284 29276 5296
rect 29227 5256 29276 5284
rect 29227 5253 29239 5256
rect 29181 5247 29239 5253
rect 29270 5244 29276 5256
rect 29328 5244 29334 5296
rect 29472 5284 29500 5324
rect 29549 5321 29561 5355
rect 29595 5352 29607 5355
rect 30466 5352 30472 5364
rect 29595 5324 30472 5352
rect 29595 5321 29607 5324
rect 29549 5315 29607 5321
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 30837 5355 30895 5361
rect 30837 5321 30849 5355
rect 30883 5321 30895 5355
rect 30837 5315 30895 5321
rect 29472 5256 29868 5284
rect 29730 5216 29736 5228
rect 27816 5188 29736 5216
rect 27157 5179 27215 5185
rect 27172 5148 27200 5179
rect 29730 5176 29736 5188
rect 29788 5176 29794 5228
rect 29840 5216 29868 5256
rect 29914 5244 29920 5296
rect 29972 5284 29978 5296
rect 30009 5287 30067 5293
rect 30009 5284 30021 5287
rect 29972 5256 30021 5284
rect 29972 5244 29978 5256
rect 30009 5253 30021 5256
rect 30055 5253 30067 5287
rect 30209 5287 30267 5293
rect 30209 5284 30221 5287
rect 30009 5247 30067 5253
rect 30208 5253 30221 5284
rect 30255 5253 30267 5287
rect 30208 5247 30267 5253
rect 30208 5216 30236 5247
rect 30852 5228 30880 5315
rect 31846 5312 31852 5364
rect 31904 5352 31910 5364
rect 32335 5355 32393 5361
rect 32335 5352 32347 5355
rect 31904 5324 32347 5352
rect 31904 5312 31910 5324
rect 32335 5321 32347 5324
rect 32381 5352 32393 5355
rect 33042 5352 33048 5364
rect 32381 5324 33048 5352
rect 32381 5321 32393 5324
rect 32335 5315 32393 5321
rect 33042 5312 33048 5324
rect 33100 5352 33106 5364
rect 33153 5355 33211 5361
rect 33153 5352 33165 5355
rect 33100 5324 33165 5352
rect 33100 5312 33106 5324
rect 33153 5321 33165 5324
rect 33199 5321 33211 5355
rect 33318 5352 33324 5364
rect 33279 5324 33324 5352
rect 33153 5315 33211 5321
rect 33318 5312 33324 5324
rect 33376 5312 33382 5364
rect 33781 5355 33839 5361
rect 33781 5321 33793 5355
rect 33827 5321 33839 5355
rect 33781 5315 33839 5321
rect 32122 5284 32128 5296
rect 32083 5256 32128 5284
rect 32122 5244 32128 5256
rect 32180 5244 32186 5296
rect 32490 5244 32496 5296
rect 32548 5284 32554 5296
rect 32953 5287 33011 5293
rect 32953 5284 32965 5287
rect 32548 5256 32965 5284
rect 32548 5244 32554 5256
rect 32953 5253 32965 5256
rect 32999 5253 33011 5287
rect 32953 5247 33011 5253
rect 29840 5188 30236 5216
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 31021 5219 31079 5225
rect 31021 5185 31033 5219
rect 31067 5185 31079 5219
rect 31021 5179 31079 5185
rect 25424 5120 27200 5148
rect 24084 5108 24090 5120
rect 22462 5080 22468 5092
rect 20496 5052 22140 5080
rect 22204 5052 22468 5080
rect 20496 5040 20502 5052
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 15528 4984 17141 5012
rect 15528 4972 15534 4984
rect 17129 4981 17141 4984
rect 17175 5012 17187 5015
rect 17218 5012 17224 5024
rect 17175 4984 17224 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18690 4972 18696 5024
rect 18748 5012 18754 5024
rect 19153 5015 19211 5021
rect 19153 5012 19165 5015
rect 18748 4984 19165 5012
rect 18748 4972 18754 4984
rect 19153 4981 19165 4984
rect 19199 4981 19211 5015
rect 19153 4975 19211 4981
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 19889 5015 19947 5021
rect 19889 5012 19901 5015
rect 19484 4984 19901 5012
rect 19484 4972 19490 4984
rect 19889 4981 19901 4984
rect 19935 4981 19947 5015
rect 19889 4975 19947 4981
rect 20809 5015 20867 5021
rect 20809 4981 20821 5015
rect 20855 5012 20867 5015
rect 21358 5012 21364 5024
rect 20855 4984 21364 5012
rect 20855 4981 20867 4984
rect 20809 4975 20867 4981
rect 21358 4972 21364 4984
rect 21416 5012 21422 5024
rect 22204 5012 22232 5052
rect 22462 5040 22468 5052
rect 22520 5040 22526 5092
rect 22646 5080 22652 5092
rect 22607 5052 22652 5080
rect 22646 5040 22652 5052
rect 22704 5040 22710 5092
rect 25314 5080 25320 5092
rect 22756 5052 25320 5080
rect 21416 4984 22232 5012
rect 21416 4972 21422 4984
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22756 5012 22784 5052
rect 25314 5040 25320 5052
rect 25372 5040 25378 5092
rect 22336 4984 22784 5012
rect 23385 5015 23443 5021
rect 22336 4972 22342 4984
rect 23385 4981 23397 5015
rect 23431 5012 23443 5015
rect 23474 5012 23480 5024
rect 23431 4984 23480 5012
rect 23431 4981 23443 4984
rect 23385 4975 23443 4981
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 24762 5012 24768 5024
rect 24723 4984 24768 5012
rect 24762 4972 24768 4984
rect 24820 4972 24826 5024
rect 25406 5012 25412 5024
rect 25367 4984 25412 5012
rect 25406 4972 25412 4984
rect 25464 4972 25470 5024
rect 26050 5012 26056 5024
rect 26011 4984 26056 5012
rect 26050 4972 26056 4984
rect 26108 4972 26114 5024
rect 26878 4972 26884 5024
rect 26936 5012 26942 5024
rect 26973 5015 27031 5021
rect 26973 5012 26985 5015
rect 26936 4984 26985 5012
rect 26936 4972 26942 4984
rect 26973 4981 26985 4984
rect 27019 4981 27031 5015
rect 26973 4975 27031 4981
rect 27062 4972 27068 5024
rect 27120 5012 27126 5024
rect 27172 5012 27200 5120
rect 27430 5108 27436 5160
rect 27488 5148 27494 5160
rect 31036 5148 31064 5179
rect 31938 5176 31944 5228
rect 31996 5216 32002 5228
rect 33796 5216 33824 5315
rect 36538 5312 36544 5364
rect 36596 5352 36602 5364
rect 36633 5355 36691 5361
rect 36633 5352 36645 5355
rect 36596 5324 36645 5352
rect 36596 5312 36602 5324
rect 36633 5321 36645 5324
rect 36679 5352 36691 5355
rect 37645 5355 37703 5361
rect 36679 5324 37320 5352
rect 36679 5321 36691 5324
rect 36633 5315 36691 5321
rect 35520 5287 35578 5293
rect 35520 5253 35532 5287
rect 35566 5284 35578 5287
rect 36262 5284 36268 5296
rect 35566 5256 36268 5284
rect 35566 5253 35578 5256
rect 35520 5247 35578 5253
rect 36262 5244 36268 5256
rect 36320 5244 36326 5296
rect 37292 5293 37320 5324
rect 37645 5321 37657 5355
rect 37691 5352 37703 5355
rect 38102 5352 38108 5364
rect 37691 5324 38108 5352
rect 37691 5321 37703 5324
rect 37645 5315 37703 5321
rect 38102 5312 38108 5324
rect 38160 5312 38166 5364
rect 37277 5287 37335 5293
rect 37277 5253 37289 5287
rect 37323 5253 37335 5287
rect 37477 5287 37535 5293
rect 37477 5284 37489 5287
rect 37277 5247 37335 5253
rect 37384 5256 37489 5284
rect 33962 5216 33968 5228
rect 31996 5188 33824 5216
rect 33923 5188 33968 5216
rect 31996 5176 32002 5188
rect 33962 5176 33968 5188
rect 34020 5176 34026 5228
rect 34609 5219 34667 5225
rect 34609 5185 34621 5219
rect 34655 5185 34667 5219
rect 34609 5179 34667 5185
rect 34624 5148 34652 5179
rect 36538 5176 36544 5228
rect 36596 5216 36602 5228
rect 37384 5216 37412 5256
rect 37477 5253 37489 5256
rect 37523 5253 37535 5287
rect 37477 5247 37535 5253
rect 36596 5188 37412 5216
rect 36596 5176 36602 5188
rect 27488 5120 31064 5148
rect 31726 5120 34652 5148
rect 27488 5108 27494 5120
rect 28445 5083 28503 5089
rect 28445 5049 28457 5083
rect 28491 5080 28503 5083
rect 28626 5080 28632 5092
rect 28491 5052 28632 5080
rect 28491 5049 28503 5052
rect 28445 5043 28503 5049
rect 28626 5040 28632 5052
rect 28684 5040 28690 5092
rect 30377 5083 30435 5089
rect 28736 5052 30328 5080
rect 28736 5012 28764 5052
rect 27120 4984 28764 5012
rect 27120 4972 27126 4984
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 29365 5015 29423 5021
rect 29365 5012 29377 5015
rect 28868 4984 29377 5012
rect 28868 4972 28874 4984
rect 29365 4981 29377 4984
rect 29411 5012 29423 5015
rect 30190 5012 30196 5024
rect 29411 4984 30196 5012
rect 29411 4981 29423 4984
rect 29365 4975 29423 4981
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 30300 5012 30328 5052
rect 30377 5049 30389 5083
rect 30423 5080 30435 5083
rect 31726 5080 31754 5120
rect 34698 5108 34704 5160
rect 34756 5148 34762 5160
rect 35253 5151 35311 5157
rect 35253 5148 35265 5151
rect 34756 5120 35265 5148
rect 34756 5108 34762 5120
rect 35253 5117 35265 5120
rect 35299 5117 35311 5151
rect 35253 5111 35311 5117
rect 30423 5052 31754 5080
rect 32493 5083 32551 5089
rect 30423 5049 30435 5052
rect 30377 5043 30435 5049
rect 32493 5049 32505 5083
rect 32539 5080 32551 5083
rect 33226 5080 33232 5092
rect 32539 5052 33232 5080
rect 32539 5049 32551 5052
rect 32493 5043 32551 5049
rect 33226 5040 33232 5052
rect 33284 5040 33290 5092
rect 34330 5040 34336 5092
rect 34388 5080 34394 5092
rect 34388 5052 35296 5080
rect 34388 5040 34394 5052
rect 31662 5012 31668 5024
rect 30300 4984 31668 5012
rect 31662 4972 31668 4984
rect 31720 4972 31726 5024
rect 31754 4972 31760 5024
rect 31812 5012 31818 5024
rect 32309 5015 32367 5021
rect 32309 5012 32321 5015
rect 31812 4984 32321 5012
rect 31812 4972 31818 4984
rect 32309 4981 32321 4984
rect 32355 5012 32367 5015
rect 32582 5012 32588 5024
rect 32355 4984 32588 5012
rect 32355 4981 32367 4984
rect 32309 4975 32367 4981
rect 32582 4972 32588 4984
rect 32640 5012 32646 5024
rect 33137 5015 33195 5021
rect 33137 5012 33149 5015
rect 32640 4984 33149 5012
rect 32640 4972 32646 4984
rect 33137 4981 33149 4984
rect 33183 4981 33195 5015
rect 34422 5012 34428 5024
rect 34383 4984 34428 5012
rect 33137 4975 33195 4981
rect 34422 4972 34428 4984
rect 34480 4972 34486 5024
rect 35268 5012 35296 5052
rect 36446 5012 36452 5024
rect 35268 4984 36452 5012
rect 36446 4972 36452 4984
rect 36504 5012 36510 5024
rect 37461 5015 37519 5021
rect 37461 5012 37473 5015
rect 36504 4984 37473 5012
rect 36504 4972 36510 4984
rect 37461 4981 37473 4984
rect 37507 4981 37519 5015
rect 37461 4975 37519 4981
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3844 4780 4752 4808
rect 3844 4768 3850 4780
rect 4724 4740 4752 4780
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 4856 4780 5273 4808
rect 4856 4768 4862 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 6914 4808 6920 4820
rect 5500 4780 6920 4808
rect 5500 4768 5506 4780
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 7616 4780 8401 4808
rect 7616 4768 7622 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 9364 4780 10241 4808
rect 9364 4768 9370 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10229 4771 10287 4777
rect 10336 4780 10701 4808
rect 5810 4740 5816 4752
rect 4724 4712 5816 4740
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 6362 4700 6368 4752
rect 6420 4740 6426 4752
rect 8570 4740 8576 4752
rect 6420 4712 8576 4740
rect 6420 4700 6426 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 9766 4740 9772 4752
rect 8956 4712 9772 4740
rect 4249 4675 4307 4681
rect 4249 4672 4261 4675
rect 3252 4644 4261 4672
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 1949 4567 2007 4573
rect 1964 4536 1992 4567
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3252 4613 3280 4644
rect 4249 4641 4261 4644
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 5994 4672 6000 4684
rect 5767 4644 6000 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 5994 4632 6000 4644
rect 6052 4672 6058 4684
rect 8956 4681 8984 4712
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 6733 4675 6791 4681
rect 6052 4644 6684 4672
rect 6052 4632 6058 4644
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3881 4607 3939 4613
rect 3881 4573 3893 4607
rect 3927 4604 3939 4607
rect 4154 4604 4160 4616
rect 3927 4576 4160 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4982 4604 4988 4616
rect 4396 4576 4988 4604
rect 4396 4564 4402 4576
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5442 4604 5448 4616
rect 5404 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 5626 4604 5632 4616
rect 5583 4576 5632 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4604 5871 4607
rect 5902 4604 5908 4616
rect 5859 4576 5908 4604
rect 5859 4573 5871 4576
rect 5813 4567 5871 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6656 4604 6684 4644
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 6779 4644 8953 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 10336 4672 10364 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 11606 4808 11612 4820
rect 11567 4780 11612 4808
rect 10689 4771 10747 4777
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 12176 4780 13461 4808
rect 12176 4752 12204 4780
rect 13449 4777 13461 4780
rect 13495 4808 13507 4811
rect 14550 4808 14556 4820
rect 13495 4780 14556 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15252 4780 15945 4808
rect 15252 4768 15258 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 25406 4808 25412 4820
rect 15933 4771 15991 4777
rect 21376 4780 25412 4808
rect 10502 4700 10508 4752
rect 10560 4700 10566 4752
rect 10962 4740 10968 4752
rect 10796 4712 10968 4740
rect 8941 4635 8999 4641
rect 9646 4644 10364 4672
rect 6822 4604 6828 4616
rect 6656 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4604 6886 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6880 4576 7021 4604
rect 6880 4564 6886 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7926 4604 7932 4616
rect 7009 4567 7067 4573
rect 7116 4576 7932 4604
rect 3786 4536 3792 4548
rect 1964 4508 3792 4536
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 4062 4536 4068 4548
rect 4023 4508 4068 4536
rect 4062 4496 4068 4508
rect 4120 4496 4126 4548
rect 7116 4536 7144 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 9214 4564 9220 4576
rect 9272 4604 9278 4616
rect 9646 4604 9674 4644
rect 10520 4613 10548 4700
rect 10796 4613 10824 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 12069 4743 12127 4749
rect 12069 4709 12081 4743
rect 12115 4740 12127 4743
rect 12158 4740 12164 4752
rect 12115 4712 12164 4740
rect 12115 4709 12127 4712
rect 12069 4703 12127 4709
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 13078 4740 13084 4752
rect 12308 4712 13084 4740
rect 12308 4700 12314 4712
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13188 4712 14228 4740
rect 13188 4672 13216 4712
rect 14090 4672 14096 4684
rect 10980 4644 13216 4672
rect 13372 4644 14096 4672
rect 9272 4576 9674 4604
rect 10396 4607 10454 4613
rect 9272 4564 9278 4576
rect 10396 4573 10408 4607
rect 10442 4604 10454 4607
rect 10506 4607 10564 4613
rect 10442 4573 10456 4604
rect 10396 4567 10456 4573
rect 10506 4573 10518 4607
rect 10552 4573 10564 4607
rect 10506 4567 10564 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 8018 4536 8024 4548
rect 4172 4508 7144 4536
rect 7979 4508 8024 4536
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 2314 4468 2320 4480
rect 1811 4440 2320 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 3234 4468 3240 4480
rect 2455 4440 3240 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 4172 4468 4200 4508
rect 8018 4496 8024 4508
rect 8076 4496 8082 4548
rect 8205 4539 8263 4545
rect 8205 4505 8217 4539
rect 8251 4536 8263 4539
rect 8662 4536 8668 4548
rect 8251 4508 8668 4536
rect 8251 4505 8263 4508
rect 8205 4499 8263 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 9950 4496 9956 4548
rect 10008 4536 10014 4548
rect 10428 4536 10456 4567
rect 10008 4508 10456 4536
rect 10008 4496 10014 4508
rect 3476 4440 4200 4468
rect 3476 4428 3482 4440
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 10980 4468 11008 4644
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11664 4576 11805 4604
rect 11664 4564 11670 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 11900 4536 11928 4567
rect 11974 4564 11980 4616
rect 12032 4604 12038 4616
rect 13372 4613 13400 4644
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 12032 4576 12173 4604
rect 12032 4564 12038 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13325 4607 13400 4613
rect 13325 4573 13337 4607
rect 13371 4576 13400 4607
rect 13371 4573 13383 4576
rect 13325 4567 13383 4573
rect 12342 4536 12348 4548
rect 11900 4508 12348 4536
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 4304 4440 11008 4468
rect 4304 4428 4310 4440
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 12250 4468 12256 4480
rect 11204 4440 12256 4468
rect 11204 4428 11210 4440
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12860 4440 13001 4468
rect 12860 4428 12866 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 13188 4468 13216 4567
rect 13446 4564 13452 4616
rect 13504 4604 13510 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13504 4576 13553 4604
rect 13504 4564 13510 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 14200 4536 14228 4712
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 21266 4740 21272 4752
rect 16724 4712 21272 4740
rect 16724 4700 16730 4712
rect 21266 4700 21272 4712
rect 21324 4700 21330 4752
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14332 4644 14565 4672
rect 14332 4632 14338 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 14568 4604 14596 4635
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 20165 4675 20223 4681
rect 20165 4672 20177 4675
rect 15620 4644 20177 4672
rect 15620 4632 15626 4644
rect 20165 4641 20177 4644
rect 20211 4641 20223 4675
rect 21376 4672 21404 4780
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 25593 4811 25651 4817
rect 25593 4777 25605 4811
rect 25639 4808 25651 4811
rect 27062 4808 27068 4820
rect 25639 4780 27068 4808
rect 25639 4777 25651 4780
rect 25593 4771 25651 4777
rect 27062 4768 27068 4780
rect 27120 4768 27126 4820
rect 28810 4808 28816 4820
rect 28771 4780 28816 4808
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 30742 4808 30748 4820
rect 28920 4780 30748 4808
rect 26050 4740 26056 4752
rect 20165 4635 20223 4641
rect 20640 4644 21404 4672
rect 22664 4712 26056 4740
rect 15102 4604 15108 4616
rect 14568 4576 15108 4604
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15286 4564 15292 4616
rect 15344 4604 15350 4616
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 15344 4576 16405 4604
rect 15344 4564 15350 4576
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 16393 4567 16451 4573
rect 16500 4576 18521 4604
rect 14798 4539 14856 4545
rect 14798 4536 14810 4539
rect 14200 4508 14810 4536
rect 14798 4505 14810 4508
rect 14844 4505 14856 4539
rect 14798 4499 14856 4505
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 16500 4536 16528 4576
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 20438 4604 20444 4616
rect 19843 4576 20444 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 20640 4613 20668 4644
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4604 22155 4607
rect 22664 4604 22692 4712
rect 26050 4700 26056 4712
rect 26108 4700 26114 4752
rect 26145 4743 26203 4749
rect 26145 4709 26157 4743
rect 26191 4709 26203 4743
rect 26145 4703 26203 4709
rect 27157 4743 27215 4749
rect 27157 4709 27169 4743
rect 27203 4740 27215 4743
rect 28920 4740 28948 4780
rect 30742 4768 30748 4780
rect 30800 4768 30806 4820
rect 31665 4811 31723 4817
rect 31665 4777 31677 4811
rect 31711 4808 31723 4811
rect 31754 4808 31760 4820
rect 31711 4780 31760 4808
rect 31711 4777 31723 4780
rect 31665 4771 31723 4777
rect 31754 4768 31760 4780
rect 31812 4768 31818 4820
rect 31849 4811 31907 4817
rect 31849 4777 31861 4811
rect 31895 4808 31907 4811
rect 32030 4808 32036 4820
rect 31895 4780 32036 4808
rect 31895 4777 31907 4780
rect 31849 4771 31907 4777
rect 32030 4768 32036 4780
rect 32088 4768 32094 4820
rect 32582 4808 32588 4820
rect 32543 4780 32588 4808
rect 32582 4768 32588 4780
rect 32640 4768 32646 4820
rect 32769 4811 32827 4817
rect 32769 4777 32781 4811
rect 32815 4808 32827 4811
rect 32815 4780 34560 4808
rect 32815 4777 32827 4780
rect 32769 4771 32827 4777
rect 27203 4712 28948 4740
rect 28997 4743 29055 4749
rect 27203 4709 27215 4712
rect 27157 4703 27215 4709
rect 28997 4709 29009 4743
rect 29043 4740 29055 4743
rect 29043 4712 31754 4740
rect 29043 4709 29055 4712
rect 28997 4703 29055 4709
rect 26160 4672 26188 4703
rect 29822 4672 29828 4684
rect 23492 4644 26188 4672
rect 28644 4644 29828 4672
rect 22830 4604 22836 4616
rect 22143 4576 22692 4604
rect 22791 4576 22836 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 15068 4508 16528 4536
rect 16577 4539 16635 4545
rect 15068 4496 15074 4508
rect 16577 4505 16589 4539
rect 16623 4536 16635 4539
rect 16666 4536 16672 4548
rect 16623 4508 16672 4536
rect 16623 4505 16635 4508
rect 16577 4499 16635 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 16758 4496 16764 4548
rect 16816 4536 16822 4548
rect 17310 4536 17316 4548
rect 16816 4508 16861 4536
rect 17271 4508 17316 4536
rect 16816 4496 16822 4508
rect 17310 4496 17316 4508
rect 17368 4496 17374 4548
rect 17497 4539 17555 4545
rect 17497 4505 17509 4539
rect 17543 4536 17555 4539
rect 18138 4536 18144 4548
rect 17543 4508 18000 4536
rect 18099 4508 18144 4536
rect 17543 4505 17555 4508
rect 17497 4499 17555 4505
rect 14274 4468 14280 4480
rect 13188 4440 14280 4468
rect 12989 4431 13047 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 17512 4468 17540 4499
rect 17678 4468 17684 4480
rect 14700 4440 17540 4468
rect 17639 4440 17684 4468
rect 14700 4428 14706 4440
rect 17678 4428 17684 4440
rect 17736 4428 17742 4480
rect 17972 4468 18000 4508
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 18325 4539 18383 4545
rect 18325 4505 18337 4539
rect 18371 4536 18383 4539
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 18371 4508 19993 4536
rect 18371 4505 18383 4508
rect 18325 4499 18383 4505
rect 19981 4505 19993 4508
rect 20027 4536 20039 4539
rect 20346 4536 20352 4548
rect 20027 4508 20352 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 18340 4468 18368 4499
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 21376 4536 21404 4567
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23492 4536 23520 4644
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 24581 4607 24639 4613
rect 23615 4576 24532 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 21376 4508 23520 4536
rect 20806 4468 20812 4480
rect 17972 4440 18368 4468
rect 20767 4440 20812 4468
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 20898 4428 20904 4480
rect 20956 4468 20962 4480
rect 21545 4471 21603 4477
rect 21545 4468 21557 4471
rect 20956 4440 21557 4468
rect 20956 4428 20962 4440
rect 21545 4437 21557 4440
rect 21591 4437 21603 4471
rect 22278 4468 22284 4480
rect 22239 4440 22284 4468
rect 21545 4431 21603 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22462 4428 22468 4480
rect 22520 4468 22526 4480
rect 23017 4471 23075 4477
rect 23017 4468 23029 4471
rect 22520 4440 23029 4468
rect 22520 4428 22526 4440
rect 23017 4437 23029 4440
rect 23063 4437 23075 4471
rect 23750 4468 23756 4480
rect 23711 4440 23756 4468
rect 23017 4431 23075 4437
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 24210 4428 24216 4480
rect 24268 4468 24274 4480
rect 24397 4471 24455 4477
rect 24397 4468 24409 4471
rect 24268 4440 24409 4468
rect 24268 4428 24274 4440
rect 24397 4437 24409 4440
rect 24443 4437 24455 4471
rect 24504 4468 24532 4576
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 24596 4536 24624 4567
rect 24670 4564 24676 4616
rect 24728 4604 24734 4616
rect 26329 4607 26387 4613
rect 26329 4604 26341 4607
rect 24728 4576 26341 4604
rect 24728 4564 24734 4576
rect 26329 4573 26341 4576
rect 26375 4573 26387 4607
rect 26878 4604 26884 4616
rect 26839 4576 26884 4604
rect 26329 4567 26387 4573
rect 26878 4564 26884 4576
rect 26936 4564 26942 4616
rect 26973 4607 27031 4613
rect 26973 4573 26985 4607
rect 27019 4604 27031 4607
rect 27154 4604 27160 4616
rect 27019 4576 27160 4604
rect 27019 4573 27031 4576
rect 26973 4567 27031 4573
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 24946 4536 24952 4548
rect 24596 4508 24952 4536
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 25314 4496 25320 4548
rect 25372 4536 25378 4548
rect 25501 4539 25559 4545
rect 25501 4536 25513 4539
rect 25372 4508 25513 4536
rect 25372 4496 25378 4508
rect 25501 4505 25513 4508
rect 25547 4505 25559 4539
rect 25501 4499 25559 4505
rect 26050 4496 26056 4548
rect 26108 4536 26114 4548
rect 26510 4536 26516 4548
rect 26108 4508 26516 4536
rect 26108 4496 26114 4508
rect 26510 4496 26516 4508
rect 26568 4496 26574 4548
rect 27062 4496 27068 4548
rect 27120 4536 27126 4548
rect 27816 4536 27844 4567
rect 28644 4545 28672 4644
rect 29822 4632 29828 4644
rect 29880 4632 29886 4684
rect 31726 4672 31754 4712
rect 32214 4700 32220 4752
rect 32272 4740 32278 4752
rect 33873 4743 33931 4749
rect 33873 4740 33885 4743
rect 32272 4712 33885 4740
rect 32272 4700 32278 4712
rect 33873 4709 33885 4712
rect 33919 4709 33931 4743
rect 34532 4740 34560 4780
rect 34606 4768 34612 4820
rect 34664 4808 34670 4820
rect 34885 4811 34943 4817
rect 34885 4808 34897 4811
rect 34664 4780 34897 4808
rect 34664 4768 34670 4780
rect 34885 4777 34897 4780
rect 34931 4777 34943 4811
rect 34885 4771 34943 4777
rect 35069 4811 35127 4817
rect 35069 4777 35081 4811
rect 35115 4808 35127 4811
rect 35342 4808 35348 4820
rect 35115 4780 35348 4808
rect 35115 4777 35127 4780
rect 35069 4771 35127 4777
rect 34900 4740 34928 4771
rect 35342 4768 35348 4780
rect 35400 4768 35406 4820
rect 35713 4811 35771 4817
rect 35713 4808 35725 4811
rect 35452 4780 35725 4808
rect 35452 4740 35480 4780
rect 35713 4777 35725 4780
rect 35759 4777 35771 4811
rect 35713 4771 35771 4777
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 35897 4811 35955 4817
rect 35897 4808 35909 4811
rect 35860 4780 35909 4808
rect 35860 4768 35866 4780
rect 35897 4777 35909 4780
rect 35943 4777 35955 4811
rect 35897 4771 35955 4777
rect 36446 4768 36452 4820
rect 36504 4808 36510 4820
rect 36633 4811 36691 4817
rect 36633 4808 36645 4811
rect 36504 4780 36645 4808
rect 36504 4768 36510 4780
rect 36633 4777 36645 4780
rect 36679 4777 36691 4811
rect 36633 4771 36691 4777
rect 36817 4811 36875 4817
rect 36817 4777 36829 4811
rect 36863 4808 36875 4811
rect 38010 4808 38016 4820
rect 36863 4780 38016 4808
rect 36863 4777 36875 4780
rect 36817 4771 36875 4777
rect 38010 4768 38016 4780
rect 38068 4768 38074 4820
rect 34532 4712 34744 4740
rect 34900 4712 35480 4740
rect 33873 4703 33931 4709
rect 33962 4672 33968 4684
rect 29932 4644 31616 4672
rect 31726 4644 33968 4672
rect 28859 4573 28917 4579
rect 27120 4508 27844 4536
rect 28629 4539 28687 4545
rect 27120 4496 27126 4508
rect 28629 4505 28641 4539
rect 28675 4505 28687 4539
rect 28859 4539 28871 4573
rect 28905 4570 28917 4573
rect 28905 4548 28939 4570
rect 29086 4564 29092 4616
rect 29144 4604 29150 4616
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29144 4576 29561 4604
rect 29144 4564 29150 4576
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4604 29791 4607
rect 29932 4604 29960 4644
rect 30760 4613 30788 4644
rect 29779 4576 29960 4604
rect 30009 4607 30067 4613
rect 29779 4573 29791 4576
rect 29733 4567 29791 4573
rect 30009 4573 30021 4607
rect 30055 4573 30067 4607
rect 30009 4567 30067 4573
rect 30745 4607 30803 4613
rect 30745 4573 30757 4607
rect 30791 4573 30803 4607
rect 31021 4607 31079 4613
rect 31021 4604 31033 4607
rect 30745 4567 30803 4573
rect 30852 4576 31033 4604
rect 28905 4539 28908 4548
rect 28859 4533 28908 4539
rect 28629 4499 28687 4505
rect 28902 4496 28908 4533
rect 28960 4496 28966 4548
rect 27617 4471 27675 4477
rect 27617 4468 27629 4471
rect 24504 4440 27629 4468
rect 24397 4431 24455 4437
rect 27617 4437 27629 4440
rect 27663 4437 27675 4471
rect 27617 4431 27675 4437
rect 28534 4428 28540 4480
rect 28592 4468 28598 4480
rect 29748 4468 29776 4567
rect 29822 4496 29828 4548
rect 29880 4536 29886 4548
rect 30024 4536 30052 4567
rect 30852 4536 30880 4576
rect 31021 4573 31033 4576
rect 31067 4573 31079 4607
rect 31021 4567 31079 4573
rect 29880 4508 30880 4536
rect 30929 4539 30987 4545
rect 29880 4496 29886 4508
rect 30929 4505 30941 4539
rect 30975 4536 30987 4539
rect 31294 4536 31300 4548
rect 30975 4508 31300 4536
rect 30975 4505 30987 4508
rect 30929 4499 30987 4505
rect 31294 4496 31300 4508
rect 31352 4536 31358 4548
rect 31481 4539 31539 4545
rect 31481 4536 31493 4539
rect 31352 4508 31493 4536
rect 31352 4496 31358 4508
rect 31481 4505 31493 4508
rect 31527 4505 31539 4539
rect 31588 4536 31616 4644
rect 33962 4632 33968 4644
rect 34020 4632 34026 4684
rect 34716 4672 34744 4712
rect 36078 4672 36084 4684
rect 34716 4644 36084 4672
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 31662 4564 31668 4616
rect 31720 4604 31726 4616
rect 31720 4576 33364 4604
rect 31720 4564 31726 4576
rect 32401 4539 32459 4545
rect 31588 4508 32260 4536
rect 31481 4499 31539 4505
rect 29914 4468 29920 4480
rect 28592 4440 29776 4468
rect 29875 4440 29920 4468
rect 28592 4428 28598 4440
rect 29914 4428 29920 4440
rect 29972 4428 29978 4480
rect 30282 4428 30288 4480
rect 30340 4468 30346 4480
rect 30561 4471 30619 4477
rect 30561 4468 30573 4471
rect 30340 4440 30573 4468
rect 30340 4428 30346 4440
rect 30561 4437 30573 4440
rect 30607 4437 30619 4471
rect 30561 4431 30619 4437
rect 31691 4471 31749 4477
rect 31691 4437 31703 4471
rect 31737 4468 31749 4471
rect 31846 4468 31852 4480
rect 31737 4440 31852 4468
rect 31737 4437 31749 4440
rect 31691 4431 31749 4437
rect 31846 4428 31852 4440
rect 31904 4428 31910 4480
rect 32232 4468 32260 4508
rect 32401 4505 32413 4539
rect 32447 4536 32459 4539
rect 32490 4536 32496 4548
rect 32447 4508 32496 4536
rect 32447 4505 32459 4508
rect 32401 4499 32459 4505
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 32617 4539 32675 4545
rect 32617 4505 32629 4539
rect 32663 4536 32675 4539
rect 33042 4536 33048 4548
rect 32663 4508 33048 4536
rect 32663 4505 32675 4508
rect 32617 4499 32675 4505
rect 33042 4496 33048 4508
rect 33100 4496 33106 4548
rect 33336 4536 33364 4576
rect 33410 4564 33416 4616
rect 33468 4604 33474 4616
rect 33468 4576 33513 4604
rect 33468 4564 33474 4576
rect 33594 4564 33600 4616
rect 33652 4604 33658 4616
rect 34057 4607 34115 4613
rect 34057 4604 34069 4607
rect 33652 4576 34069 4604
rect 33652 4564 33658 4576
rect 34057 4573 34069 4576
rect 34103 4573 34115 4607
rect 36538 4604 36544 4616
rect 34057 4567 34115 4573
rect 34624 4576 36544 4604
rect 34624 4536 34652 4576
rect 36538 4564 36544 4576
rect 36596 4564 36602 4616
rect 37642 4564 37648 4616
rect 37700 4604 37706 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 37700 4576 37841 4604
rect 37700 4564 37706 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 33336 4508 34652 4536
rect 34701 4539 34759 4545
rect 34701 4505 34713 4539
rect 34747 4536 34759 4539
rect 34790 4536 34796 4548
rect 34747 4508 34796 4536
rect 34747 4505 34759 4508
rect 34701 4499 34759 4505
rect 34790 4496 34796 4508
rect 34848 4496 34854 4548
rect 34882 4496 34888 4548
rect 34940 4545 34946 4548
rect 34940 4539 34959 4545
rect 34947 4536 34959 4539
rect 35529 4539 35587 4545
rect 34947 4508 35020 4536
rect 34947 4505 34959 4508
rect 34940 4499 34959 4505
rect 34940 4496 34946 4499
rect 32306 4468 32312 4480
rect 32232 4440 32312 4468
rect 32306 4428 32312 4440
rect 32364 4428 32370 4480
rect 33226 4468 33232 4480
rect 33187 4440 33232 4468
rect 33226 4428 33232 4440
rect 33284 4428 33290 4480
rect 33410 4428 33416 4480
rect 33468 4468 33474 4480
rect 34238 4468 34244 4480
rect 33468 4440 34244 4468
rect 33468 4428 33474 4440
rect 34238 4428 34244 4440
rect 34296 4428 34302 4480
rect 34992 4468 35020 4508
rect 35529 4505 35541 4539
rect 35575 4536 35587 4539
rect 36078 4536 36084 4548
rect 35575 4508 36084 4536
rect 35575 4505 35587 4508
rect 35529 4499 35587 4505
rect 36078 4496 36084 4508
rect 36136 4496 36142 4548
rect 36170 4496 36176 4548
rect 36228 4536 36234 4548
rect 36449 4539 36507 4545
rect 36449 4536 36461 4539
rect 36228 4508 36461 4536
rect 36228 4496 36234 4508
rect 36449 4505 36461 4508
rect 36495 4505 36507 4539
rect 36556 4536 36584 4564
rect 36649 4539 36707 4545
rect 36649 4536 36661 4539
rect 36556 4508 36661 4536
rect 36449 4499 36507 4505
rect 36649 4505 36661 4508
rect 36695 4505 36707 4539
rect 36649 4499 36707 4505
rect 35729 4471 35787 4477
rect 35729 4468 35741 4471
rect 34992 4440 35741 4468
rect 35729 4437 35741 4440
rect 35775 4437 35787 4471
rect 35729 4431 35787 4437
rect 37918 4428 37924 4480
rect 37976 4468 37982 4480
rect 38013 4471 38071 4477
rect 38013 4468 38025 4471
rect 37976 4440 38025 4468
rect 37976 4428 37982 4440
rect 38013 4437 38025 4440
rect 38059 4437 38071 4471
rect 38013 4431 38071 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2869 4267 2927 4273
rect 2372 4236 2774 4264
rect 2372 4224 2378 4236
rect 2746 4196 2774 4236
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 3418 4264 3424 4276
rect 2915 4236 3424 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 4246 4264 4252 4276
rect 3559 4236 4252 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4706 4264 4712 4276
rect 4448 4236 4712 4264
rect 2746 4168 2912 4196
rect 2884 4140 2912 4168
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 1872 3992 1900 4091
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3602 4128 3608 4140
rect 3099 4100 3608 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 3878 4128 3884 4140
rect 3743 4100 3884 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4338 4128 4344 4140
rect 4299 4100 4344 4128
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4448 4137 4476 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 7374 4264 7380 4276
rect 6564 4236 7380 4264
rect 6564 4196 6592 4236
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 8018 4264 8024 4276
rect 7515 4236 8024 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 11698 4264 11704 4276
rect 8720 4236 11704 4264
rect 8720 4224 8726 4236
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 13078 4264 13084 4276
rect 12032 4236 13084 4264
rect 12032 4224 12038 4236
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 13633 4267 13691 4273
rect 13633 4233 13645 4267
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 5460 4168 6592 4196
rect 5460 4140 5488 4168
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4531 4128 4568 4132
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4531 4100 4721 4128
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 4531 4060 4559 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 4709 4091 4767 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5442 4128 5448 4140
rect 5403 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 5810 4128 5816 4140
rect 5592 4100 5637 4128
rect 5771 4100 5816 4128
rect 5592 4088 5598 4100
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 6564 4137 6592 4168
rect 7006 4156 7012 4208
rect 7064 4196 7070 4208
rect 7064 4168 8138 4196
rect 7064 4156 7070 4168
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6730 4128 6736 4140
rect 6687 4100 6736 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7432 4100 7665 4128
rect 7432 4088 7438 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 8018 4128 8024 4140
rect 7791 4100 7880 4128
rect 7979 4100 8024 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 7852 4072 7880 4100
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8110 4128 8138 4168
rect 8570 4156 8576 4208
rect 8628 4196 8634 4208
rect 9582 4196 9588 4208
rect 8628 4168 9588 4196
rect 8628 4156 8634 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 9674 4156 9680 4208
rect 9732 4156 9738 4208
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 10468 4168 11529 4196
rect 10468 4156 10474 4168
rect 11517 4165 11529 4168
rect 11563 4165 11575 4199
rect 12802 4196 12808 4208
rect 11517 4159 11575 4165
rect 11624 4168 11928 4196
rect 12763 4168 12808 4196
rect 9692 4128 9720 4156
rect 11624 4128 11652 4168
rect 8110 4100 9720 4128
rect 9784 4100 11652 4128
rect 2372 4032 4559 4060
rect 4617 4063 4675 4069
rect 2372 4020 2378 4032
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 5350 4060 5356 4072
rect 4663 4032 5356 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 7558 4060 7564 4072
rect 5552 4032 7564 4060
rect 3418 3992 3424 4004
rect 1872 3964 3424 3992
rect 3418 3952 3424 3964
rect 3476 3952 3482 4004
rect 3694 3952 3700 4004
rect 3752 3992 3758 4004
rect 5442 3992 5448 4004
rect 3752 3964 5448 3992
rect 3752 3952 3758 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 5552 3924 5580 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 9784 4069 9812 4100
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 11900 4128 11928 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 12989 4199 13047 4205
rect 12989 4165 13001 4199
rect 13035 4196 13047 4199
rect 13262 4196 13268 4208
rect 13035 4168 13268 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 13648 4196 13676 4227
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 15194 4264 15200 4276
rect 14332 4236 15200 4264
rect 14332 4224 14338 4236
rect 15194 4224 15200 4236
rect 15252 4264 15258 4276
rect 15252 4236 15608 4264
rect 15252 4224 15258 4236
rect 14642 4196 14648 4208
rect 13648 4168 14648 4196
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 14918 4196 14924 4208
rect 14752 4168 14924 4196
rect 13170 4128 13176 4140
rect 11756 4100 11801 4128
rect 11900 4100 12756 4128
rect 13131 4100 13176 4128
rect 11756 4088 11762 4100
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8260 4032 8493 4060
rect 8260 4020 8266 4032
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 8527 4032 9781 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 10008 4032 10057 4060
rect 10008 4020 10014 4032
rect 10045 4029 10057 4032
rect 10091 4060 10103 4063
rect 11606 4060 11612 4072
rect 10091 4032 11612 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 12728 4060 12756 4100
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 14182 4128 14188 4140
rect 13863 4100 14188 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 14332 4100 14473 4128
rect 14332 4088 14338 4100
rect 14461 4097 14473 4100
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 14752 4128 14780 4168
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 14599 4100 14780 4128
rect 14829 4131 14887 4137
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 14829 4097 14841 4131
rect 14875 4128 14887 4131
rect 14875 4100 15424 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 12728 4032 14412 4060
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 11974 3992 11980 4004
rect 5684 3964 11980 3992
rect 5684 3952 5690 3964
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 1719 3896 5580 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 5994 3924 6000 3936
rect 5776 3896 6000 3924
rect 5776 3884 5782 3896
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 7984 3896 8029 3924
rect 7984 3884 7990 3896
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8711 3927 8769 3933
rect 8711 3924 8723 3927
rect 8628 3896 8723 3924
rect 8628 3884 8634 3896
rect 8711 3893 8723 3896
rect 8757 3893 8769 3927
rect 8711 3887 8769 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 11146 3924 11152 3936
rect 8996 3896 11152 3924
rect 8996 3884 9002 3896
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11882 3924 11888 3936
rect 11388 3896 11888 3924
rect 11388 3884 11394 3896
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 14274 3924 14280 3936
rect 14235 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 14384 3924 14412 4032
rect 14660 4032 14749 4060
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 14660 3992 14688 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 15286 4060 15292 4072
rect 15247 4032 15292 4060
rect 14737 4023 14795 4029
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 14608 3964 14688 3992
rect 14608 3952 14614 3964
rect 15304 3924 15332 4020
rect 15396 3992 15424 4100
rect 15580 4069 15608 4236
rect 16298 4224 16304 4276
rect 16356 4264 16362 4276
rect 18046 4264 18052 4276
rect 16356 4236 18052 4264
rect 16356 4224 16362 4236
rect 18046 4224 18052 4236
rect 18104 4264 18110 4276
rect 20438 4264 20444 4276
rect 18104 4236 20024 4264
rect 20399 4236 20444 4264
rect 18104 4224 18110 4236
rect 19610 4196 19616 4208
rect 19168 4168 19616 4196
rect 19168 4140 19196 4168
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 19996 4196 20024 4236
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 22554 4224 22560 4276
rect 22612 4264 22618 4276
rect 27341 4267 27399 4273
rect 22612 4236 26464 4264
rect 22612 4224 22618 4236
rect 19996 4168 20668 4196
rect 16850 4088 16856 4140
rect 16908 4128 16914 4140
rect 16908 4100 16953 4128
rect 16908 4088 16914 4100
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 18874 4137 18880 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17276 4100 17325 4128
rect 17276 4088 17282 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 18868 4128 18880 4137
rect 18835 4100 18880 4128
rect 17313 4091 17371 4097
rect 18868 4091 18880 4100
rect 18874 4088 18880 4091
rect 18932 4088 18938 4140
rect 19150 4088 19156 4140
rect 19208 4088 19214 4140
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 20162 4128 20168 4140
rect 19300 4100 20168 4128
rect 19300 4088 19306 4100
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20640 4137 20668 4168
rect 21266 4156 21272 4208
rect 21324 4196 21330 4208
rect 24026 4196 24032 4208
rect 21324 4168 24032 4196
rect 21324 4156 21330 4168
rect 24026 4156 24032 4168
rect 24084 4156 24090 4208
rect 24486 4156 24492 4208
rect 24544 4196 24550 4208
rect 26436 4196 26464 4236
rect 27341 4233 27353 4267
rect 27387 4264 27399 4267
rect 27430 4264 27436 4276
rect 27387 4236 27436 4264
rect 27387 4233 27399 4236
rect 27341 4227 27399 4233
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 29454 4264 29460 4276
rect 27540 4236 29460 4264
rect 27540 4196 27568 4236
rect 29454 4224 29460 4236
rect 29512 4224 29518 4276
rect 29549 4267 29607 4273
rect 29549 4233 29561 4267
rect 29595 4264 29607 4267
rect 29914 4264 29920 4276
rect 29595 4236 29920 4264
rect 29595 4233 29607 4236
rect 29549 4227 29607 4233
rect 29914 4224 29920 4236
rect 29972 4224 29978 4276
rect 30190 4224 30196 4276
rect 30248 4264 30254 4276
rect 33226 4264 33232 4276
rect 30248 4236 33232 4264
rect 30248 4224 30254 4236
rect 33226 4224 33232 4236
rect 33284 4224 33290 4276
rect 34606 4224 34612 4276
rect 34664 4264 34670 4276
rect 35545 4267 35603 4273
rect 35545 4264 35557 4267
rect 34664 4236 35557 4264
rect 34664 4224 34670 4236
rect 35545 4233 35557 4236
rect 35591 4233 35603 4267
rect 35545 4227 35603 4233
rect 29086 4196 29092 4208
rect 24544 4168 25176 4196
rect 26436 4168 27568 4196
rect 28644 4168 29092 4196
rect 24544 4156 24550 4168
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4097 20683 4131
rect 20625 4091 20683 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20990 4128 20996 4140
rect 20772 4100 20817 4128
rect 20951 4100 20996 4128
rect 20772 4088 20778 4100
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 22370 4128 22376 4140
rect 22327 4100 22376 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22548 4131 22606 4137
rect 22548 4097 22560 4131
rect 22594 4128 22606 4131
rect 23474 4128 23480 4140
rect 22594 4100 23480 4128
rect 22594 4097 22606 4100
rect 22548 4091 22606 4097
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 24394 4128 24400 4140
rect 24355 4100 24400 4128
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24670 4128 24676 4140
rect 24627 4100 24676 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 24820 4100 25053 4128
rect 24820 4088 24826 4100
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25148 4128 25176 4168
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 25148 4100 25237 4128
rect 25041 4091 25099 4097
rect 25225 4097 25237 4100
rect 25271 4097 25283 4131
rect 25225 4091 25283 4097
rect 25409 4131 25467 4137
rect 25409 4097 25421 4131
rect 25455 4128 25467 4131
rect 25682 4128 25688 4140
rect 25455 4100 25688 4128
rect 25455 4097 25467 4100
rect 25409 4091 25467 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 25866 4088 25872 4140
rect 25924 4128 25930 4140
rect 26237 4131 26295 4137
rect 26237 4128 26249 4131
rect 25924 4100 26249 4128
rect 25924 4088 25930 4100
rect 26237 4097 26249 4100
rect 26283 4097 26295 4131
rect 26418 4128 26424 4140
rect 26379 4100 26424 4128
rect 26237 4091 26295 4097
rect 26418 4088 26424 4100
rect 26476 4088 26482 4140
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26936 4100 26985 4128
rect 26936 4088 26942 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4128 27215 4131
rect 27338 4128 27344 4140
rect 27203 4100 27344 4128
rect 27203 4097 27215 4100
rect 27157 4091 27215 4097
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 28166 4128 28172 4140
rect 28127 4100 28172 4128
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 28436 4131 28494 4137
rect 28436 4097 28448 4131
rect 28482 4128 28494 4131
rect 28644 4128 28672 4168
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 29822 4156 29828 4208
rect 29880 4196 29886 4208
rect 35345 4199 35403 4205
rect 29880 4168 31754 4196
rect 29880 4156 29886 4168
rect 28482 4100 28672 4128
rect 28482 4097 28494 4100
rect 28436 4091 28494 4097
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 30006 4128 30012 4140
rect 28868 4100 30012 4128
rect 28868 4088 28874 4100
rect 30006 4088 30012 4100
rect 30064 4088 30070 4140
rect 30282 4137 30288 4140
rect 30276 4128 30288 4137
rect 30243 4100 30288 4128
rect 30276 4091 30288 4100
rect 30282 4088 30288 4091
rect 30340 4088 30346 4140
rect 31726 4128 31754 4168
rect 32232 4168 32628 4196
rect 32232 4128 32260 4168
rect 31726 4100 32260 4128
rect 32306 4088 32312 4140
rect 32364 4128 32370 4140
rect 32490 4128 32496 4140
rect 32364 4100 32409 4128
rect 32451 4100 32496 4128
rect 32364 4088 32370 4100
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 32600 4137 32628 4168
rect 35345 4165 35357 4199
rect 35391 4196 35403 4199
rect 35434 4196 35440 4208
rect 35391 4168 35440 4196
rect 35391 4165 35403 4168
rect 35345 4159 35403 4165
rect 35434 4156 35440 4168
rect 35492 4156 35498 4208
rect 32585 4131 32643 4137
rect 32585 4097 32597 4131
rect 32631 4128 32643 4131
rect 33318 4128 33324 4140
rect 32631 4100 33324 4128
rect 32631 4097 32643 4100
rect 32585 4091 32643 4097
rect 33318 4088 33324 4100
rect 33376 4088 33382 4140
rect 33772 4131 33830 4137
rect 33772 4097 33784 4131
rect 33818 4128 33830 4131
rect 34514 4128 34520 4140
rect 33818 4100 34520 4128
rect 33818 4097 33830 4100
rect 33772 4091 33830 4097
rect 34514 4088 34520 4100
rect 34572 4088 34578 4140
rect 36449 4131 36507 4137
rect 36449 4097 36461 4131
rect 36495 4128 36507 4131
rect 36722 4128 36728 4140
rect 36495 4100 36728 4128
rect 36495 4097 36507 4100
rect 36449 4091 36507 4097
rect 36722 4088 36728 4100
rect 36780 4088 36786 4140
rect 37274 4128 37280 4140
rect 37235 4100 37280 4128
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16206 4060 16212 4072
rect 15611 4032 16212 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4060 17647 4063
rect 18230 4060 18236 4072
rect 17635 4032 18236 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18598 4060 18604 4072
rect 18559 4032 18604 4060
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 19760 4032 20913 4060
rect 19760 4020 19766 4032
rect 20901 4029 20913 4032
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4060 24271 4063
rect 24780 4060 24808 4088
rect 24259 4032 24808 4060
rect 26053 4063 26111 4069
rect 24259 4029 24271 4032
rect 24213 4023 24271 4029
rect 26053 4029 26065 4063
rect 26099 4060 26111 4063
rect 26510 4060 26516 4072
rect 26099 4032 26516 4060
rect 26099 4029 26111 4032
rect 26053 4023 26111 4029
rect 26510 4020 26516 4032
rect 26568 4060 26574 4072
rect 26896 4060 26924 4088
rect 26568 4032 26924 4060
rect 26568 4020 26574 4032
rect 32122 4020 32128 4072
rect 32180 4060 32186 4072
rect 33505 4063 33563 4069
rect 33505 4060 33517 4063
rect 32180 4032 33517 4060
rect 32180 4020 32186 4032
rect 33505 4029 33517 4032
rect 33551 4029 33563 4063
rect 37182 4060 37188 4072
rect 33505 4023 33563 4029
rect 35728 4032 37188 4060
rect 15654 3992 15660 4004
rect 15396 3964 15660 3992
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 33410 3992 33416 4004
rect 23348 3964 27016 3992
rect 23348 3952 23354 3964
rect 16666 3924 16672 3936
rect 14384 3896 15332 3924
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 19794 3924 19800 3936
rect 17092 3896 19800 3924
rect 17092 3884 17098 3896
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20162 3924 20168 3936
rect 20027 3896 20168 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 23474 3884 23480 3936
rect 23532 3924 23538 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23532 3896 23673 3924
rect 23532 3884 23538 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 24946 3884 24952 3936
rect 25004 3924 25010 3936
rect 26878 3924 26884 3936
rect 25004 3896 26884 3924
rect 25004 3884 25010 3896
rect 26878 3884 26884 3896
rect 26936 3884 26942 3936
rect 26988 3924 27016 3964
rect 30944 3964 33416 3992
rect 30944 3924 30972 3964
rect 33410 3952 33416 3964
rect 33468 3952 33474 4004
rect 26988 3896 30972 3924
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 31389 3927 31447 3933
rect 31389 3924 31401 3927
rect 31352 3896 31401 3924
rect 31352 3884 31358 3896
rect 31389 3893 31401 3896
rect 31435 3893 31447 3927
rect 31389 3887 31447 3893
rect 31478 3884 31484 3936
rect 31536 3924 31542 3936
rect 32125 3927 32183 3933
rect 32125 3924 32137 3927
rect 31536 3896 32137 3924
rect 31536 3884 31542 3896
rect 32125 3893 32137 3896
rect 32171 3893 32183 3927
rect 33520 3924 33548 4023
rect 35728 4001 35756 4032
rect 37182 4020 37188 4032
rect 37240 4020 37246 4072
rect 35713 3995 35771 4001
rect 35713 3961 35725 3995
rect 35759 3961 35771 3995
rect 35713 3955 35771 3961
rect 36633 3995 36691 4001
rect 36633 3961 36645 3995
rect 36679 3992 36691 3995
rect 38654 3992 38660 4004
rect 36679 3964 38660 3992
rect 36679 3961 36691 3964
rect 36633 3955 36691 3961
rect 38654 3952 38660 3964
rect 38712 3952 38718 4004
rect 34698 3924 34704 3936
rect 33520 3896 34704 3924
rect 32125 3887 32183 3893
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 34885 3927 34943 3933
rect 34885 3924 34897 3927
rect 34848 3896 34897 3924
rect 34848 3884 34854 3896
rect 34885 3893 34897 3896
rect 34931 3893 34943 3927
rect 34885 3887 34943 3893
rect 35434 3884 35440 3936
rect 35492 3924 35498 3936
rect 35529 3927 35587 3933
rect 35529 3924 35541 3927
rect 35492 3896 35541 3924
rect 35492 3884 35498 3896
rect 35529 3893 35541 3896
rect 35575 3893 35587 3927
rect 35529 3887 35587 3893
rect 37182 3884 37188 3936
rect 37240 3924 37246 3936
rect 37461 3927 37519 3933
rect 37461 3924 37473 3927
rect 37240 3896 37473 3924
rect 37240 3884 37246 3896
rect 37461 3893 37473 3896
rect 37507 3893 37519 3927
rect 37461 3887 37519 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3326 3720 3332 3732
rect 2332 3692 3332 3720
rect 2332 3661 2360 3692
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 6788 3692 7021 3720
rect 6788 3680 6794 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 7009 3683 7067 3689
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 12250 3720 12256 3732
rect 7340 3692 12256 3720
rect 7340 3680 7346 3692
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 15378 3720 15384 3732
rect 13320 3692 15384 3720
rect 13320 3680 13326 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17221 3723 17279 3729
rect 17221 3720 17233 3723
rect 17000 3692 17233 3720
rect 17000 3680 17006 3692
rect 17221 3689 17233 3692
rect 17267 3689 17279 3723
rect 17221 3683 17279 3689
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3621 2375 3655
rect 2317 3615 2375 3621
rect 5169 3655 5227 3661
rect 5169 3621 5181 3655
rect 5215 3652 5227 3655
rect 5534 3652 5540 3664
rect 5215 3624 5540 3652
rect 5215 3621 5227 3624
rect 5169 3615 5227 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 8021 3655 8079 3661
rect 8021 3621 8033 3655
rect 8067 3652 8079 3655
rect 8110 3652 8116 3664
rect 8067 3624 8116 3652
rect 8067 3621 8079 3624
rect 8021 3615 8079 3621
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 8938 3652 8944 3664
rect 8168 3624 8944 3652
rect 8168 3612 8174 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 9968 3624 10333 3652
rect 3694 3584 3700 3596
rect 1688 3556 3700 3584
rect 1688 3525 1716 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 8570 3584 8576 3596
rect 7432 3556 8576 3584
rect 7432 3544 7438 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 1820 3488 1865 3516
rect 1820 3476 1826 3488
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 3234 3516 3240 3528
rect 2004 3488 2049 3516
rect 3195 3488 3240 3516
rect 2004 3476 2010 3488
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4614 3516 4620 3528
rect 3835 3488 4620 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4614 3476 4620 3488
rect 4672 3516 4678 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 4672 3488 5641 3516
rect 4672 3476 4678 3488
rect 5629 3485 5641 3488
rect 5675 3516 5687 3519
rect 6730 3516 6736 3528
rect 5675 3488 6736 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6730 3476 6736 3488
rect 6788 3516 6794 3528
rect 7760 3525 7788 3556
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 8904 3556 9076 3584
rect 8904 3544 8910 3556
rect 7745 3519 7803 3525
rect 6788 3488 7697 3516
rect 6788 3476 6794 3488
rect 4034 3451 4092 3457
rect 4034 3448 4046 3451
rect 3068 3420 4046 3448
rect 3068 3389 3096 3420
rect 4034 3417 4046 3420
rect 4080 3417 4092 3451
rect 4034 3411 4092 3417
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 5874 3451 5932 3457
rect 5874 3448 5886 3451
rect 5776 3420 5886 3448
rect 5776 3408 5782 3420
rect 5874 3417 5886 3420
rect 5920 3417 5932 3451
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 5874 3411 5932 3417
rect 7484 3420 7573 3448
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 7282 3380 7288 3392
rect 3936 3352 7288 3380
rect 3936 3340 3942 3352
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 7484 3380 7512 3420
rect 7561 3417 7573 3420
rect 7607 3417 7619 3451
rect 7669 3448 7697 3488
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8110 3516 8116 3528
rect 7892 3488 7937 3516
rect 8071 3488 8116 3516
rect 7892 3476 7898 3488
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 9048 3516 9076 3556
rect 9968 3516 9996 3624
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 12345 3655 12403 3661
rect 12345 3652 12357 3655
rect 12124 3624 12357 3652
rect 12124 3612 12130 3624
rect 12345 3621 12357 3624
rect 12391 3621 12403 3655
rect 12345 3615 12403 3621
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15838 3584 15844 3596
rect 15160 3556 15844 3584
rect 15160 3544 15166 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 17236 3584 17264 3683
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17368 3692 17877 3720
rect 17368 3680 17374 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 18782 3720 18788 3732
rect 18380 3692 18788 3720
rect 18380 3680 18386 3692
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 18966 3680 18972 3732
rect 19024 3720 19030 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 19024 3692 19257 3720
rect 19024 3680 19030 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 19702 3720 19708 3732
rect 19392 3692 19708 3720
rect 19392 3680 19398 3692
rect 19702 3680 19708 3692
rect 19760 3720 19766 3732
rect 20349 3723 20407 3729
rect 20349 3720 20361 3723
rect 19760 3692 20361 3720
rect 19760 3680 19766 3692
rect 20349 3689 20361 3692
rect 20395 3689 20407 3723
rect 22370 3720 22376 3732
rect 20349 3683 20407 3689
rect 20916 3692 22376 3720
rect 17589 3655 17647 3661
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 17635 3624 18460 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 17236 3556 18184 3584
rect 11238 3525 11244 3528
rect 9048 3488 9996 3516
rect 10965 3519 11023 3525
rect 8941 3479 8999 3485
rect 10965 3485 10977 3519
rect 11011 3485 11023 3519
rect 11232 3516 11244 3525
rect 11199 3488 11244 3516
rect 10965 3479 11023 3485
rect 11232 3479 11244 3488
rect 8956 3448 8984 3479
rect 7669 3420 8984 3448
rect 7561 3411 7619 3417
rect 7432 3352 7512 3380
rect 8956 3380 8984 3420
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9186 3451 9244 3457
rect 9186 3448 9198 3451
rect 9088 3420 9198 3448
rect 9088 3408 9094 3420
rect 9186 3417 9198 3420
rect 9232 3417 9244 3451
rect 9186 3411 9244 3417
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 10980 3448 11008 3479
rect 11238 3476 11244 3479
rect 11296 3476 11302 3528
rect 12434 3516 12440 3528
rect 11348 3488 12440 3516
rect 11348 3448 11376 3488
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 12986 3516 12992 3528
rect 12584 3488 12992 3516
rect 12584 3476 12590 3488
rect 12986 3476 12992 3488
rect 13044 3516 13050 3528
rect 13262 3516 13268 3528
rect 13044 3488 13268 3516
rect 13044 3476 13050 3488
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14260 3519 14318 3525
rect 14260 3516 14272 3519
rect 14148 3488 14272 3516
rect 14148 3476 14154 3488
rect 14260 3485 14272 3488
rect 14306 3485 14318 3519
rect 14260 3479 14318 3485
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14642 3516 14648 3528
rect 14424 3488 14469 3516
rect 14603 3488 14648 3516
rect 14424 3476 14430 3488
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 18156 3525 18184 3556
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 18288 3556 18337 3584
rect 18288 3544 18294 3556
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 18325 3547 18383 3553
rect 18432 3584 18460 3624
rect 18598 3612 18604 3664
rect 18656 3652 18662 3664
rect 18656 3624 20668 3652
rect 18656 3612 18662 3624
rect 20346 3584 20352 3596
rect 18432 3556 19334 3584
rect 18432 3525 18460 3556
rect 16097 3519 16155 3525
rect 16097 3516 16109 3519
rect 15252 3488 16109 3516
rect 15252 3476 15258 3488
rect 16097 3485 16109 3488
rect 16143 3485 16155 3519
rect 16097 3479 16155 3485
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 9364 3420 10456 3448
rect 10980 3420 11376 3448
rect 9364 3408 9370 3420
rect 9582 3380 9588 3392
rect 8956 3352 9588 3380
rect 7432 3340 7438 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10318 3380 10324 3392
rect 9732 3352 10324 3380
rect 9732 3340 9738 3352
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10428 3380 10456 3420
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 11572 3420 12817 3448
rect 11572 3408 11578 3420
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 13170 3448 13176 3460
rect 13131 3420 13176 3448
rect 12805 3411 12863 3417
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 13924 3420 14228 3448
rect 13924 3380 13952 3420
rect 14090 3380 14096 3392
rect 10428 3352 13952 3380
rect 14051 3352 14096 3380
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14200 3380 14228 3420
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 15105 3451 15163 3457
rect 15105 3448 15117 3451
rect 14884 3420 15117 3448
rect 14884 3408 14890 3420
rect 15105 3417 15117 3420
rect 15151 3417 15163 3451
rect 15105 3411 15163 3417
rect 15289 3451 15347 3457
rect 15289 3417 15301 3451
rect 15335 3448 15347 3451
rect 15378 3448 15384 3460
rect 15335 3420 15384 3448
rect 15335 3417 15347 3420
rect 15289 3411 15347 3417
rect 15378 3408 15384 3420
rect 15436 3408 15442 3460
rect 15473 3383 15531 3389
rect 15473 3380 15485 3383
rect 14200 3352 15485 3380
rect 15473 3349 15485 3352
rect 15519 3349 15531 3383
rect 15473 3343 15531 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 18064 3380 18092 3479
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 19058 3448 19064 3460
rect 18288 3420 19064 3448
rect 18288 3408 18294 3420
rect 19058 3408 19064 3420
rect 19116 3408 19122 3460
rect 19306 3448 19334 3556
rect 19444 3556 20352 3584
rect 19444 3525 19472 3556
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20640 3584 20668 3624
rect 20916 3593 20944 3692
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 25685 3723 25743 3729
rect 25685 3689 25697 3723
rect 25731 3720 25743 3723
rect 26234 3720 26240 3732
rect 25731 3692 26240 3720
rect 25731 3689 25743 3692
rect 25685 3683 25743 3689
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 27893 3723 27951 3729
rect 27893 3689 27905 3723
rect 27939 3720 27951 3723
rect 28994 3720 29000 3732
rect 27939 3692 29000 3720
rect 27939 3689 27951 3692
rect 27893 3683 27951 3689
rect 28994 3680 29000 3692
rect 29052 3680 29058 3732
rect 32401 3723 32459 3729
rect 32401 3689 32413 3723
rect 32447 3720 32459 3723
rect 32490 3720 32496 3732
rect 32447 3692 32496 3720
rect 32447 3689 32459 3692
rect 32401 3683 32459 3689
rect 32490 3680 32496 3692
rect 32548 3680 32554 3732
rect 33962 3720 33968 3732
rect 33923 3692 33968 3720
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 34146 3720 34152 3732
rect 34107 3692 34152 3720
rect 34146 3680 34152 3692
rect 34204 3680 34210 3732
rect 35434 3720 35440 3732
rect 34716 3692 35440 3720
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 23750 3652 23756 3664
rect 23164 3624 23756 3652
rect 23164 3612 23170 3624
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 25593 3655 25651 3661
rect 23860 3624 25544 3652
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20640 3556 20913 3584
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19944 3488 20085 3516
rect 19944 3476 19950 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20441 3519 20499 3525
rect 20211 3488 20300 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 19518 3448 19524 3460
rect 19306 3420 19524 3448
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 19904 3448 19932 3476
rect 19812 3420 19932 3448
rect 19812 3380 19840 3420
rect 17460 3352 19840 3380
rect 19889 3383 19947 3389
rect 17460 3340 17466 3352
rect 19889 3349 19901 3383
rect 19935 3380 19947 3383
rect 20162 3380 20168 3392
rect 19935 3352 20168 3380
rect 19935 3349 19947 3352
rect 19889 3343 19947 3349
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 20272 3380 20300 3488
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 20530 3516 20536 3528
rect 20487 3488 20536 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20640 3448 20668 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 20901 3547 20959 3553
rect 23382 3544 23388 3596
rect 23440 3584 23446 3596
rect 23860 3584 23888 3624
rect 24765 3587 24823 3593
rect 24765 3584 24777 3587
rect 23440 3556 23888 3584
rect 24136 3556 24777 3584
rect 23440 3544 23446 3556
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20990 3516 20996 3528
rect 20772 3488 20996 3516
rect 20772 3476 20778 3488
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 22833 3479 22891 3485
rect 20806 3448 20812 3460
rect 20640 3420 20812 3448
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 21174 3457 21180 3460
rect 21168 3411 21180 3457
rect 21232 3448 21238 3460
rect 22848 3448 22876 3479
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23845 3519 23903 3525
rect 23247 3488 23796 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23474 3448 23480 3460
rect 21232 3420 21268 3448
rect 22848 3420 23480 3448
rect 21174 3408 21180 3411
rect 21232 3408 21238 3420
rect 23474 3408 23480 3420
rect 23532 3408 23538 3460
rect 21450 3380 21456 3392
rect 20272 3352 21456 3380
rect 21450 3340 21456 3352
rect 21508 3380 21514 3392
rect 22281 3383 22339 3389
rect 22281 3380 22293 3383
rect 21508 3352 22293 3380
rect 21508 3340 21514 3352
rect 22281 3349 22293 3352
rect 22327 3349 22339 3383
rect 22281 3343 22339 3349
rect 23290 3340 23296 3392
rect 23348 3380 23354 3392
rect 23661 3383 23719 3389
rect 23661 3380 23673 3383
rect 23348 3352 23673 3380
rect 23348 3340 23354 3352
rect 23661 3349 23673 3352
rect 23707 3349 23719 3383
rect 23768 3380 23796 3488
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 24136 3516 24164 3556
rect 24765 3553 24777 3556
rect 24811 3553 24823 3587
rect 25516 3584 25544 3624
rect 25593 3621 25605 3655
rect 25639 3652 25651 3655
rect 26510 3652 26516 3664
rect 25639 3624 26516 3652
rect 25639 3621 25651 3624
rect 25593 3615 25651 3621
rect 26510 3612 26516 3624
rect 26568 3612 26574 3664
rect 27801 3655 27859 3661
rect 27801 3621 27813 3655
rect 27847 3652 27859 3655
rect 28902 3652 28908 3664
rect 27847 3624 28908 3652
rect 27847 3621 27859 3624
rect 27801 3615 27859 3621
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 33980 3652 34008 3680
rect 34330 3652 34336 3664
rect 33980 3624 34336 3652
rect 34330 3612 34336 3624
rect 34388 3652 34394 3664
rect 34716 3652 34744 3692
rect 35434 3680 35440 3692
rect 35492 3720 35498 3732
rect 36078 3720 36084 3732
rect 35492 3692 35940 3720
rect 36039 3692 36084 3720
rect 35492 3680 35498 3692
rect 34388 3624 34744 3652
rect 35912 3652 35940 3692
rect 36078 3680 36084 3692
rect 36136 3680 36142 3732
rect 36725 3723 36783 3729
rect 36725 3720 36737 3723
rect 36188 3692 36737 3720
rect 36188 3652 36216 3692
rect 36725 3689 36737 3692
rect 36771 3689 36783 3723
rect 36906 3720 36912 3732
rect 36867 3692 36912 3720
rect 36725 3683 36783 3689
rect 36906 3680 36912 3692
rect 36964 3680 36970 3732
rect 35912 3624 36216 3652
rect 34388 3612 34394 3624
rect 36446 3612 36452 3664
rect 36504 3652 36510 3664
rect 37553 3655 37611 3661
rect 37553 3652 37565 3655
rect 36504 3624 37565 3652
rect 36504 3612 36510 3624
rect 37553 3621 37565 3624
rect 37599 3621 37611 3655
rect 37553 3615 37611 3621
rect 25866 3584 25872 3596
rect 25516 3556 25872 3584
rect 24765 3547 24823 3553
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 26050 3544 26056 3596
rect 26108 3584 26114 3596
rect 26145 3587 26203 3593
rect 26145 3584 26157 3587
rect 26108 3556 26157 3584
rect 26108 3544 26114 3556
rect 26145 3553 26157 3556
rect 26191 3553 26203 3587
rect 26145 3547 26203 3553
rect 27246 3544 27252 3596
rect 27304 3584 27310 3596
rect 27433 3587 27491 3593
rect 27433 3584 27445 3587
rect 27304 3556 27445 3584
rect 27304 3544 27310 3556
rect 27433 3553 27445 3556
rect 27479 3553 27491 3587
rect 27433 3547 27491 3553
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28718 3584 28724 3596
rect 27764 3556 28724 3584
rect 27764 3544 27770 3556
rect 28718 3544 28724 3556
rect 28776 3544 28782 3596
rect 29822 3584 29828 3596
rect 28920 3556 29828 3584
rect 23891 3488 24164 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24268 3488 24409 3516
rect 24268 3476 24274 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 26602 3516 26608 3528
rect 24627 3488 26608 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 26602 3476 26608 3488
rect 26660 3476 26666 3528
rect 26878 3476 26884 3528
rect 26936 3516 26942 3528
rect 26936 3488 27752 3516
rect 26936 3476 26942 3488
rect 25225 3451 25283 3457
rect 25225 3417 25237 3451
rect 25271 3448 25283 3451
rect 27614 3448 27620 3460
rect 25271 3420 27620 3448
rect 25271 3417 25283 3420
rect 25225 3411 25283 3417
rect 27614 3408 27620 3420
rect 27672 3408 27678 3460
rect 27724 3448 27752 3488
rect 27798 3476 27804 3528
rect 27856 3516 27862 3528
rect 28258 3516 28264 3528
rect 27856 3488 28264 3516
rect 27856 3476 27862 3488
rect 28258 3476 28264 3488
rect 28316 3476 28322 3528
rect 28626 3516 28632 3528
rect 28587 3488 28632 3516
rect 28626 3476 28632 3488
rect 28684 3476 28690 3528
rect 28920 3525 28948 3556
rect 29822 3544 29828 3556
rect 29880 3544 29886 3596
rect 30006 3544 30012 3596
rect 30064 3584 30070 3596
rect 31021 3587 31079 3593
rect 31021 3584 31033 3587
rect 30064 3556 31033 3584
rect 30064 3544 30070 3556
rect 31021 3553 31033 3556
rect 31067 3553 31079 3587
rect 31021 3547 31079 3553
rect 28905 3519 28963 3525
rect 28905 3485 28917 3519
rect 28951 3485 28963 3519
rect 28905 3479 28963 3485
rect 29549 3519 29607 3525
rect 29549 3485 29561 3519
rect 29595 3516 29607 3519
rect 29730 3516 29736 3528
rect 29595 3488 29736 3516
rect 29595 3485 29607 3488
rect 29549 3479 29607 3485
rect 29730 3476 29736 3488
rect 29788 3516 29794 3528
rect 30190 3516 30196 3528
rect 29788 3488 30196 3516
rect 29788 3476 29794 3488
rect 30190 3476 30196 3488
rect 30248 3476 30254 3528
rect 31036 3516 31064 3547
rect 32858 3544 32864 3596
rect 32916 3584 32922 3596
rect 34698 3584 34704 3596
rect 32916 3556 34040 3584
rect 34659 3556 34704 3584
rect 32916 3544 32922 3556
rect 32122 3516 32128 3528
rect 31036 3488 32128 3516
rect 32122 3476 32128 3488
rect 32180 3476 32186 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 32364 3488 33057 3516
rect 32364 3476 32370 3488
rect 33045 3485 33057 3488
rect 33091 3485 33103 3519
rect 33318 3516 33324 3528
rect 33279 3488 33324 3516
rect 33045 3479 33103 3485
rect 33318 3476 33324 3488
rect 33376 3476 33382 3528
rect 34012 3516 34040 3556
rect 34698 3544 34704 3556
rect 34756 3544 34762 3596
rect 34606 3516 34612 3528
rect 34012 3491 34612 3516
rect 34011 3488 34612 3491
rect 34011 3485 34069 3488
rect 31110 3448 31116 3460
rect 27724 3420 31116 3448
rect 31110 3408 31116 3420
rect 31168 3408 31174 3460
rect 31288 3451 31346 3457
rect 31288 3417 31300 3451
rect 31334 3448 31346 3451
rect 31478 3448 31484 3460
rect 31334 3420 31484 3448
rect 31334 3417 31346 3420
rect 31288 3411 31346 3417
rect 31478 3408 31484 3420
rect 31536 3408 31542 3460
rect 33229 3451 33287 3457
rect 33229 3417 33241 3451
rect 33275 3448 33287 3451
rect 33502 3448 33508 3460
rect 33275 3420 33508 3448
rect 33275 3417 33287 3420
rect 33229 3411 33287 3417
rect 33502 3408 33508 3420
rect 33560 3448 33566 3460
rect 33781 3451 33839 3457
rect 33781 3448 33793 3451
rect 33560 3420 33793 3448
rect 33560 3408 33566 3420
rect 33781 3417 33793 3420
rect 33827 3417 33839 3451
rect 34011 3451 34023 3485
rect 34057 3451 34069 3485
rect 34606 3476 34612 3488
rect 34664 3476 34670 3528
rect 37366 3516 37372 3528
rect 37327 3488 37372 3516
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 34011 3445 34069 3451
rect 34968 3451 35026 3457
rect 33781 3411 33839 3417
rect 34968 3417 34980 3451
rect 35014 3448 35026 3451
rect 35618 3448 35624 3460
rect 35014 3420 35624 3448
rect 35014 3417 35026 3420
rect 34968 3411 35026 3417
rect 35618 3408 35624 3420
rect 35676 3408 35682 3460
rect 36078 3408 36084 3460
rect 36136 3448 36142 3460
rect 36541 3451 36599 3457
rect 36541 3448 36553 3451
rect 36136 3420 36553 3448
rect 36136 3408 36142 3420
rect 36541 3417 36553 3420
rect 36587 3417 36599 3451
rect 36541 3411 36599 3417
rect 24026 3380 24032 3392
rect 23768 3352 24032 3380
rect 23661 3343 23719 3349
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 24118 3340 24124 3392
rect 24176 3380 24182 3392
rect 26605 3383 26663 3389
rect 26605 3380 26617 3383
rect 24176 3352 26617 3380
rect 24176 3340 24182 3352
rect 26605 3349 26617 3352
rect 26651 3349 26663 3383
rect 26605 3343 26663 3349
rect 27246 3340 27252 3392
rect 27304 3380 27310 3392
rect 27890 3380 27896 3392
rect 27304 3352 27896 3380
rect 27304 3340 27310 3352
rect 27890 3340 27896 3352
rect 27948 3340 27954 3392
rect 28442 3380 28448 3392
rect 28403 3352 28448 3380
rect 28442 3340 28448 3352
rect 28500 3340 28506 3392
rect 28813 3383 28871 3389
rect 28813 3349 28825 3383
rect 28859 3380 28871 3383
rect 29086 3380 29092 3392
rect 28859 3352 29092 3380
rect 28859 3349 28871 3352
rect 28813 3343 28871 3349
rect 29086 3340 29092 3352
rect 29144 3340 29150 3392
rect 32858 3380 32864 3392
rect 32819 3352 32864 3380
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 36722 3340 36728 3392
rect 36780 3389 36786 3392
rect 36780 3383 36799 3389
rect 36787 3349 36799 3383
rect 36780 3343 36799 3349
rect 36780 3340 36786 3343
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3142 3176 3148 3188
rect 3007 3148 3148 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3973 3179 4031 3185
rect 3973 3176 3985 3179
rect 3292 3148 3985 3176
rect 3292 3136 3298 3148
rect 3973 3145 3985 3148
rect 4019 3145 4031 3179
rect 3973 3139 4031 3145
rect 4062 3136 4068 3188
rect 4120 3136 4126 3188
rect 4982 3176 4988 3188
rect 4632 3148 4988 3176
rect 3602 3108 3608 3120
rect 3563 3080 3608 3108
rect 3602 3068 3608 3080
rect 3660 3068 3666 3120
rect 3789 3111 3847 3117
rect 3789 3077 3801 3111
rect 3835 3108 3847 3111
rect 4080 3108 4108 3136
rect 3835 3080 4108 3108
rect 3835 3077 3847 3080
rect 3789 3071 3847 3077
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4632 3049 4660 3148
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 6880 3148 7043 3176
rect 6880 3136 6886 3148
rect 5445 3111 5503 3117
rect 4724 3080 5304 3108
rect 4724 3049 4752 3080
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5166 3040 5172 3052
rect 5031 3012 5172 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5276 3040 5304 3080
rect 5445 3077 5457 3111
rect 5491 3108 5503 3111
rect 6362 3108 6368 3120
rect 5491 3080 6368 3108
rect 5491 3077 5503 3080
rect 5445 3071 5503 3077
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 7015 3117 7043 3148
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 8076 3148 8125 3176
rect 8076 3136 8082 3148
rect 8113 3145 8125 3148
rect 8159 3176 8171 3179
rect 8478 3176 8484 3188
rect 8159 3148 8484 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8628 3148 14596 3176
rect 8628 3136 8634 3148
rect 6989 3111 7047 3117
rect 6989 3077 7001 3111
rect 7035 3077 7047 3111
rect 6989 3071 7047 3077
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7248 3080 10916 3108
rect 7248 3068 7254 3080
rect 5534 3040 5540 3052
rect 5276 3012 5540 3040
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 6086 3040 6092 3052
rect 5675 3012 6092 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 7558 3040 7564 3052
rect 6840 3012 7564 3040
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6840 2972 6868 3012
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 6604 2944 6868 2972
rect 8772 2972 8800 3003
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9122 3040 9128 3052
rect 8904 3012 8949 3040
rect 9083 3012 9128 3040
rect 8904 3000 8910 3012
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9841 3043 9899 3049
rect 9841 3040 9853 3043
rect 9692 3012 9853 3040
rect 9490 2972 9496 2984
rect 8772 2944 9496 2972
rect 6604 2932 6610 2944
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9692 2972 9720 3012
rect 9841 3009 9853 3012
rect 9887 3009 9899 3043
rect 9841 3003 9899 3009
rect 9600 2944 9720 2972
rect 10888 2972 10916 3080
rect 12544 3080 14412 3108
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 11974 3040 11980 3052
rect 11839 3012 11980 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 11514 2972 11520 2984
rect 10888 2944 11376 2972
rect 11475 2944 11520 2972
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 4433 2907 4491 2913
rect 4433 2904 4445 2907
rect 3660 2876 4445 2904
rect 3660 2864 3666 2876
rect 4433 2873 4445 2876
rect 4479 2873 4491 2907
rect 4433 2867 4491 2873
rect 4816 2876 6776 2904
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2836 1731 2839
rect 4816 2836 4844 2876
rect 1719 2808 4844 2836
rect 4893 2839 4951 2845
rect 1719 2805 1731 2808
rect 1673 2799 1731 2805
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 5626 2836 5632 2848
rect 4939 2808 5632 2836
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 6748 2836 6776 2876
rect 8110 2836 8116 2848
rect 6748 2808 8116 2836
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8570 2836 8576 2848
rect 8531 2808 8576 2836
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 9214 2836 9220 2848
rect 9079 2808 9220 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 9214 2796 9220 2808
rect 9272 2836 9278 2848
rect 9398 2836 9404 2848
rect 9272 2808 9404 2836
rect 9272 2796 9278 2808
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 9600 2836 9628 2944
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10836 2876 10977 2904
rect 10836 2864 10842 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 11348 2904 11376 2944
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 12084 2972 12112 3003
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12544 3049 12572 3080
rect 14384 3049 14412 3080
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12492 3012 12541 3040
rect 12492 3000 12498 3012
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12785 3043 12843 3049
rect 12785 3040 12797 3043
rect 12529 3003 12587 3009
rect 12636 3012 12797 3040
rect 11900 2944 12112 2972
rect 11900 2904 11928 2944
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12636 2972 12664 3012
rect 12785 3009 12797 3012
rect 12831 3009 12843 3043
rect 12785 3003 12843 3009
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14568 3040 14596 3148
rect 14918 3136 14924 3188
rect 14976 3176 14982 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 14976 3148 15761 3176
rect 14976 3136 14982 3148
rect 15749 3145 15761 3148
rect 15795 3145 15807 3179
rect 15749 3139 15807 3145
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 19426 3176 19432 3188
rect 16908 3148 19432 3176
rect 16908 3136 16914 3148
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 20806 3176 20812 3188
rect 20088 3148 20812 3176
rect 15838 3068 15844 3120
rect 15896 3108 15902 3120
rect 15896 3080 17080 3108
rect 15896 3068 15902 3080
rect 14625 3043 14683 3049
rect 14625 3040 14637 3043
rect 14568 3012 14637 3040
rect 14369 3003 14427 3009
rect 14625 3009 14637 3012
rect 14671 3009 14683 3043
rect 14625 3003 14683 3009
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 16022 3040 16028 3052
rect 15436 3012 16028 3040
rect 15436 3000 15442 3012
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 17052 3049 17080 3080
rect 18046 3068 18052 3120
rect 18104 3108 18110 3120
rect 18104 3080 18552 3108
rect 18104 3068 18110 3080
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17293 3043 17351 3049
rect 17293 3040 17305 3043
rect 17037 3003 17095 3009
rect 17144 3012 17305 3040
rect 17144 2972 17172 3012
rect 17293 3009 17305 3012
rect 17339 3009 17351 3043
rect 18524 3040 18552 3080
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18524 3012 19073 3040
rect 17293 3003 17351 3009
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19242 3040 19248 3052
rect 19199 3012 19248 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 19383 3043 19441 3049
rect 19383 3009 19395 3043
rect 19429 3040 19441 3043
rect 19794 3040 19800 3052
rect 19429 3012 19800 3040
rect 19429 3009 19441 3012
rect 19383 3003 19441 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3040 19947 3043
rect 20088 3040 20116 3148
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 23017 3179 23075 3185
rect 23017 3145 23029 3179
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 23845 3179 23903 3185
rect 23845 3145 23857 3179
rect 23891 3176 23903 3179
rect 24302 3176 24308 3188
rect 23891 3148 24308 3176
rect 23891 3145 23903 3148
rect 23845 3139 23903 3145
rect 20346 3068 20352 3120
rect 20404 3108 20410 3120
rect 23032 3108 23060 3139
rect 24302 3136 24308 3148
rect 24360 3136 24366 3188
rect 25317 3179 25375 3185
rect 25317 3145 25329 3179
rect 25363 3176 25375 3179
rect 25590 3176 25596 3188
rect 25363 3148 25596 3176
rect 25363 3145 25375 3148
rect 25317 3139 25375 3145
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 26142 3176 26148 3188
rect 26103 3148 26148 3176
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 29086 3176 29092 3188
rect 29047 3148 29092 3176
rect 29086 3136 29092 3148
rect 29144 3176 29150 3188
rect 29144 3148 29592 3176
rect 29144 3136 29150 3148
rect 20404 3080 23060 3108
rect 20404 3068 20410 3080
rect 24026 3068 24032 3120
rect 24084 3108 24090 3120
rect 28166 3108 28172 3120
rect 24084 3080 24532 3108
rect 24084 3068 24090 3080
rect 19935 3012 20116 3040
rect 20156 3043 20214 3049
rect 19935 3009 19947 3012
rect 19889 3003 19947 3009
rect 20156 3009 20168 3043
rect 20202 3040 20214 3043
rect 20438 3040 20444 3052
rect 20202 3012 20444 3040
rect 20202 3009 20214 3012
rect 20156 3003 20214 3009
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 20530 3000 20536 3052
rect 20588 3040 20594 3052
rect 21450 3040 21456 3052
rect 20588 3012 21456 3040
rect 20588 3000 20594 3012
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21560 3012 22017 3040
rect 12308 2944 12664 2972
rect 15396 2944 17172 2972
rect 12308 2932 12314 2944
rect 11348 2876 11928 2904
rect 11977 2907 12035 2913
rect 10965 2867 11023 2873
rect 11977 2873 11989 2907
rect 12023 2904 12035 2907
rect 12158 2904 12164 2916
rect 12023 2876 12164 2904
rect 12023 2873 12035 2876
rect 11977 2867 12035 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 13909 2907 13967 2913
rect 13909 2873 13921 2907
rect 13955 2904 13967 2907
rect 14366 2904 14372 2916
rect 13955 2876 14372 2904
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 14366 2864 14372 2876
rect 14424 2864 14430 2916
rect 11790 2836 11796 2848
rect 9600 2808 11796 2836
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 15396 2836 15424 2944
rect 21082 2932 21088 2984
rect 21140 2972 21146 2984
rect 21560 2972 21588 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 23382 3040 23388 3052
rect 22879 3012 23388 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 21140 2944 21588 2972
rect 21821 2975 21879 2981
rect 21140 2932 21146 2944
rect 21821 2941 21833 2975
rect 21867 2972 21879 2975
rect 22756 2972 22784 3003
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 23658 3040 23664 3052
rect 23619 3012 23664 3040
rect 23658 3000 23664 3012
rect 23716 3000 23722 3052
rect 24504 3049 24532 3080
rect 27724 3080 28172 3108
rect 24489 3043 24547 3049
rect 24489 3009 24501 3043
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 24762 3000 24768 3052
rect 24820 3040 24826 3052
rect 24949 3043 25007 3049
rect 24949 3040 24961 3043
rect 24820 3012 24961 3040
rect 24820 3000 24826 3012
rect 24949 3009 24961 3012
rect 24995 3009 25007 3043
rect 24949 3003 25007 3009
rect 25133 3043 25191 3049
rect 25133 3009 25145 3043
rect 25179 3040 25191 3043
rect 25222 3040 25228 3052
rect 25179 3012 25228 3040
rect 25179 3009 25191 3012
rect 25133 3003 25191 3009
rect 23474 2972 23480 2984
rect 21867 2944 23480 2972
rect 21867 2941 21879 2944
rect 21821 2935 21879 2941
rect 23474 2932 23480 2944
rect 23532 2972 23538 2984
rect 24210 2972 24216 2984
rect 23532 2944 24216 2972
rect 23532 2932 23538 2944
rect 24210 2932 24216 2944
rect 24268 2932 24274 2984
rect 24964 2972 24992 3003
rect 25222 3000 25228 3012
rect 25280 3000 25286 3052
rect 25958 3040 25964 3052
rect 25919 3012 25964 3040
rect 25958 3000 25964 3012
rect 26016 3000 26022 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 27724 3049 27752 3080
rect 28166 3068 28172 3080
rect 28224 3068 28230 3120
rect 29564 3117 29592 3148
rect 30006 3136 30012 3188
rect 30064 3176 30070 3188
rect 31297 3179 31355 3185
rect 31297 3176 31309 3179
rect 30064 3148 31309 3176
rect 30064 3136 30070 3148
rect 31297 3145 31309 3148
rect 31343 3145 31355 3179
rect 33502 3176 33508 3188
rect 33463 3148 33508 3176
rect 31297 3139 31355 3145
rect 33502 3136 33508 3148
rect 33560 3136 33566 3188
rect 34606 3136 34612 3188
rect 34664 3176 34670 3188
rect 34993 3179 35051 3185
rect 34993 3176 35005 3179
rect 34664 3148 35005 3176
rect 34664 3136 34670 3148
rect 34993 3145 35005 3148
rect 35039 3145 35051 3179
rect 34993 3139 35051 3145
rect 35161 3179 35219 3185
rect 35161 3145 35173 3179
rect 35207 3176 35219 3179
rect 36173 3179 36231 3185
rect 35207 3148 36124 3176
rect 35207 3145 35219 3148
rect 35161 3139 35219 3145
rect 29549 3111 29607 3117
rect 29549 3077 29561 3111
rect 29595 3077 29607 3111
rect 29749 3111 29807 3117
rect 29749 3108 29761 3111
rect 29549 3071 29607 3077
rect 29656 3080 29761 3108
rect 27709 3043 27767 3049
rect 27709 3009 27721 3043
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 27798 3000 27804 3052
rect 27856 3000 27862 3052
rect 27976 3043 28034 3049
rect 27976 3009 27988 3043
rect 28022 3040 28034 3043
rect 28442 3040 28448 3052
rect 28022 3012 28448 3040
rect 28022 3009 28034 3012
rect 27976 3003 28034 3009
rect 28442 3000 28448 3012
rect 28500 3000 28506 3052
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 29656 3040 29684 3080
rect 29749 3077 29761 3080
rect 29795 3077 29807 3111
rect 32214 3108 32220 3120
rect 29749 3071 29807 3077
rect 30392 3080 32220 3108
rect 30392 3049 30420 3080
rect 32214 3068 32220 3080
rect 32272 3068 32278 3120
rect 32392 3111 32450 3117
rect 32392 3077 32404 3111
rect 32438 3108 32450 3111
rect 32858 3108 32864 3120
rect 32438 3080 32864 3108
rect 32438 3077 32450 3080
rect 32392 3071 32450 3077
rect 32858 3068 32864 3080
rect 32916 3068 32922 3120
rect 34790 3108 34796 3120
rect 34751 3080 34796 3108
rect 34790 3068 34796 3080
rect 34848 3068 34854 3120
rect 28960 3012 29684 3040
rect 30377 3043 30435 3049
rect 28960 3000 28966 3012
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 31113 3043 31171 3049
rect 31113 3009 31125 3043
rect 31159 3040 31171 3043
rect 31938 3040 31944 3052
rect 31159 3012 31944 3040
rect 31159 3009 31171 3012
rect 31113 3003 31171 3009
rect 31938 3000 31944 3012
rect 31996 3000 32002 3052
rect 32122 3040 32128 3052
rect 32083 3012 32128 3040
rect 32122 3000 32128 3012
rect 32180 3000 32186 3052
rect 33594 3040 33600 3052
rect 32232 3012 33600 3040
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 24964 2944 25789 2972
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 25866 2932 25872 2984
rect 25924 2972 25930 2984
rect 27816 2972 27844 3000
rect 25924 2944 27844 2972
rect 25924 2932 25930 2944
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 31386 2972 31392 2984
rect 28776 2944 31392 2972
rect 28776 2932 28782 2944
rect 31386 2932 31392 2944
rect 31444 2932 31450 2984
rect 32232 2972 32260 3012
rect 33594 3000 33600 3012
rect 33652 3000 33658 3052
rect 33686 3000 33692 3052
rect 33744 3040 33750 3052
rect 33965 3043 34023 3049
rect 33965 3040 33977 3043
rect 33744 3012 33977 3040
rect 33744 3000 33750 3012
rect 33965 3009 33977 3012
rect 34011 3009 34023 3043
rect 35008 3040 35036 3139
rect 35805 3111 35863 3117
rect 35805 3077 35817 3111
rect 35851 3108 35863 3111
rect 35894 3108 35900 3120
rect 35851 3080 35900 3108
rect 35851 3077 35863 3080
rect 35805 3071 35863 3077
rect 35894 3068 35900 3080
rect 35952 3068 35958 3120
rect 36005 3111 36063 3117
rect 36005 3077 36017 3111
rect 36051 3077 36063 3111
rect 36096 3108 36124 3148
rect 36173 3145 36185 3179
rect 36219 3176 36231 3179
rect 36630 3176 36636 3188
rect 36219 3148 36636 3176
rect 36219 3145 36231 3148
rect 36173 3139 36231 3145
rect 36630 3136 36636 3148
rect 36688 3136 36694 3188
rect 36814 3108 36820 3120
rect 36096 3080 36820 3108
rect 36005 3071 36063 3077
rect 36020 3040 36048 3071
rect 36814 3068 36820 3080
rect 36872 3068 36878 3120
rect 36722 3040 36728 3052
rect 35008 3012 36728 3040
rect 33965 3003 34023 3009
rect 36722 3000 36728 3012
rect 36780 3000 36786 3052
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37458 3040 37464 3052
rect 37323 3012 37464 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 31726 2944 32260 2972
rect 18322 2864 18328 2916
rect 18380 2904 18386 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 18380 2876 18429 2904
rect 18380 2864 18386 2876
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 22189 2907 22247 2913
rect 22189 2904 22201 2907
rect 18417 2867 18475 2873
rect 20824 2876 22201 2904
rect 12492 2808 15424 2836
rect 12492 2796 12498 2808
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 18230 2836 18236 2848
rect 16172 2808 18236 2836
rect 16172 2796 16178 2808
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 18874 2836 18880 2848
rect 18835 2808 18880 2836
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 19334 2836 19340 2848
rect 19295 2808 19340 2836
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19610 2796 19616 2848
rect 19668 2836 19674 2848
rect 20824 2836 20852 2876
rect 22189 2873 22201 2876
rect 22235 2873 22247 2907
rect 22189 2867 22247 2873
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 22796 2876 24440 2904
rect 22796 2864 22802 2876
rect 19668 2808 20852 2836
rect 19668 2796 19674 2808
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 21269 2839 21327 2845
rect 21269 2836 21281 2839
rect 21048 2808 21281 2836
rect 21048 2796 21054 2808
rect 21269 2805 21281 2808
rect 21315 2805 21327 2839
rect 21269 2799 21327 2805
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 22278 2836 22284 2848
rect 21692 2808 22284 2836
rect 21692 2796 21698 2808
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 24302 2836 24308 2848
rect 24263 2808 24308 2836
rect 24302 2796 24308 2808
rect 24360 2796 24366 2848
rect 24412 2836 24440 2876
rect 25314 2864 25320 2916
rect 25372 2904 25378 2916
rect 27157 2907 27215 2913
rect 27157 2904 27169 2907
rect 25372 2876 27169 2904
rect 25372 2864 25378 2876
rect 27157 2873 27169 2876
rect 27203 2873 27215 2907
rect 27706 2904 27712 2916
rect 27157 2867 27215 2873
rect 27264 2876 27712 2904
rect 27264 2836 27292 2876
rect 27706 2864 27712 2876
rect 27764 2864 27770 2916
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 29917 2907 29975 2913
rect 29144 2876 29868 2904
rect 29144 2864 29150 2876
rect 24412 2808 27292 2836
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 28994 2836 29000 2848
rect 27672 2808 29000 2836
rect 27672 2796 27678 2808
rect 28994 2796 29000 2808
rect 29052 2796 29058 2848
rect 29730 2836 29736 2848
rect 29691 2808 29736 2836
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 29840 2836 29868 2876
rect 29917 2873 29929 2907
rect 29963 2904 29975 2907
rect 31726 2904 31754 2944
rect 29963 2876 31754 2904
rect 29963 2873 29975 2876
rect 29917 2867 29975 2873
rect 35710 2864 35716 2916
rect 35768 2904 35774 2916
rect 37461 2907 37519 2913
rect 37461 2904 37473 2907
rect 35768 2876 37473 2904
rect 35768 2864 35774 2876
rect 37461 2873 37473 2876
rect 37507 2873 37519 2907
rect 37461 2867 37519 2873
rect 30561 2839 30619 2845
rect 30561 2836 30573 2839
rect 29840 2808 30573 2836
rect 30561 2805 30573 2808
rect 30607 2805 30619 2839
rect 30561 2799 30619 2805
rect 32766 2796 32772 2848
rect 32824 2836 32830 2848
rect 34149 2839 34207 2845
rect 34149 2836 34161 2839
rect 32824 2808 34161 2836
rect 32824 2796 32830 2808
rect 34149 2805 34161 2808
rect 34195 2805 34207 2839
rect 34149 2799 34207 2805
rect 34330 2796 34336 2848
rect 34388 2836 34394 2848
rect 34977 2839 35035 2845
rect 34977 2836 34989 2839
rect 34388 2808 34989 2836
rect 34388 2796 34394 2808
rect 34977 2805 34989 2808
rect 35023 2836 35035 2839
rect 35989 2839 36047 2845
rect 35989 2836 36001 2839
rect 35023 2808 36001 2836
rect 35023 2805 35035 2808
rect 34977 2799 35035 2805
rect 35989 2805 36001 2808
rect 36035 2805 36047 2839
rect 35989 2799 36047 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 5534 2632 5540 2644
rect 3016 2604 5540 2632
rect 3016 2592 3022 2604
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 5718 2632 5724 2644
rect 5675 2604 5724 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 9030 2632 9036 2644
rect 8251 2604 9036 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10410 2632 10416 2644
rect 9999 2604 10416 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 12434 2632 12440 2644
rect 11655 2604 12440 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 13814 2632 13820 2644
rect 12544 2604 13820 2632
rect 2682 2524 2688 2576
rect 2740 2564 2746 2576
rect 4985 2567 5043 2573
rect 2740 2536 4844 2564
rect 2740 2524 2746 2536
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3878 2496 3884 2508
rect 3283 2468 3884 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4816 2496 4844 2536
rect 4985 2533 4997 2567
rect 5031 2564 5043 2567
rect 12250 2564 12256 2576
rect 5031 2536 12256 2564
rect 5031 2533 5043 2536
rect 4985 2527 5043 2533
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 12544 2564 12572 2604
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 15194 2632 15200 2644
rect 14507 2604 15200 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15930 2592 15936 2644
rect 15988 2632 15994 2644
rect 17678 2632 17684 2644
rect 15988 2604 17684 2632
rect 15988 2592 15994 2604
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 18138 2632 18144 2644
rect 18095 2604 18144 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 18782 2632 18788 2644
rect 18656 2604 18788 2632
rect 18656 2592 18662 2604
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 19613 2635 19671 2641
rect 19613 2601 19625 2635
rect 19659 2632 19671 2635
rect 20070 2632 20076 2644
rect 19659 2604 20076 2632
rect 19659 2601 19671 2604
rect 19613 2595 19671 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20533 2635 20591 2641
rect 20533 2601 20545 2635
rect 20579 2632 20591 2635
rect 20622 2632 20628 2644
rect 20579 2604 20628 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 20732 2604 27292 2632
rect 15289 2567 15347 2573
rect 12406 2536 12572 2564
rect 12820 2536 15240 2564
rect 6822 2496 6828 2508
rect 4816 2468 6828 2496
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 6932 2468 7757 2496
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6932 2437 6960 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 7745 2459 7803 2465
rect 8404 2468 9321 2496
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 6917 2391 6975 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 8404 2437 8432 2468
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 9456 2468 10425 2496
rect 9456 2456 9462 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 12406 2496 12434 2536
rect 10413 2459 10471 2465
rect 11808 2468 12434 2496
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8628 2400 8953 2428
rect 8628 2388 8634 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 10008 2400 10149 2428
rect 10008 2388 10014 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 10229 2391 10287 2397
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 624 2332 1869 2360
rect 624 2320 630 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2041 2363 2099 2369
rect 2041 2329 2053 2363
rect 2087 2360 2099 2363
rect 7282 2360 7288 2372
rect 2087 2332 7288 2360
rect 2087 2329 2099 2332
rect 2041 2323 2099 2329
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7561 2363 7619 2369
rect 7561 2329 7573 2363
rect 7607 2360 7619 2363
rect 8478 2360 8484 2372
rect 7607 2332 8484 2360
rect 7607 2329 7619 2332
rect 7561 2323 7619 2329
rect 8478 2320 8484 2332
rect 8536 2360 8542 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8536 2332 9137 2360
rect 8536 2320 8542 2332
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 10244 2360 10272 2391
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 11808 2437 11836 2468
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12820 2428 12848 2536
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 15010 2496 15016 2508
rect 13872 2468 15016 2496
rect 13872 2456 13878 2468
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 15212 2496 15240 2536
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 17218 2564 17224 2576
rect 15335 2536 17224 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2564 17371 2567
rect 17494 2564 17500 2576
rect 17359 2536 17500 2564
rect 17359 2533 17371 2536
rect 17313 2527 17371 2533
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2564 18567 2567
rect 19334 2564 19340 2576
rect 18555 2536 19340 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 15562 2496 15568 2508
rect 15212 2468 15568 2496
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 16666 2496 16672 2508
rect 15856 2468 16672 2496
rect 12483 2400 12848 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 15856 2437 15884 2468
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 18782 2456 18788 2508
rect 18840 2496 18846 2508
rect 20732 2496 20760 2604
rect 24578 2524 24584 2576
rect 24636 2564 24642 2576
rect 25777 2567 25835 2573
rect 25777 2564 25789 2567
rect 24636 2536 25789 2564
rect 24636 2524 24642 2536
rect 25777 2533 25789 2536
rect 25823 2533 25835 2567
rect 25777 2527 25835 2533
rect 23290 2496 23296 2508
rect 18840 2468 20760 2496
rect 21008 2468 23296 2496
rect 18840 2456 18846 2468
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 13044 2400 13093 2428
rect 13044 2388 13050 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 10870 2360 10876 2372
rect 10244 2332 10876 2360
rect 9125 2323 9183 2329
rect 10870 2320 10876 2332
rect 10928 2320 10934 2372
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 14090 2360 14096 2372
rect 12943 2332 14096 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 14090 2320 14096 2332
rect 14148 2320 14154 2372
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3200 2264 3985 2292
rect 3200 2252 3206 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 12250 2292 12256 2304
rect 12211 2264 12256 2292
rect 3973 2255 4031 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 13262 2292 13268 2304
rect 13223 2264 13268 2292
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 14660 2292 14688 2391
rect 15120 2360 15148 2391
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 16264 2400 17141 2428
rect 16264 2388 16270 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18233 2431 18291 2437
rect 18233 2428 18245 2431
rect 18104 2400 18245 2428
rect 18104 2388 18110 2400
rect 18233 2397 18245 2400
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 18322 2388 18328 2440
rect 18380 2428 18386 2440
rect 18598 2428 18604 2440
rect 18380 2400 18425 2428
rect 18559 2400 18604 2428
rect 18380 2388 18386 2400
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18932 2400 19257 2428
rect 18932 2388 18938 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 19518 2428 19524 2440
rect 19475 2400 19524 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 20162 2428 20168 2440
rect 20123 2400 20168 2428
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 21008 2437 21036 2468
rect 23290 2456 23296 2468
rect 23348 2456 23354 2508
rect 24762 2496 24768 2508
rect 24723 2468 24768 2496
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2496 25191 2499
rect 27062 2496 27068 2508
rect 25179 2468 27068 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 27062 2456 27068 2468
rect 27120 2456 27126 2508
rect 27264 2505 27292 2604
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 29052 2604 30481 2632
rect 29052 2592 29058 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 30469 2595 30527 2601
rect 32030 2592 32036 2644
rect 32088 2632 32094 2644
rect 33781 2635 33839 2641
rect 33781 2632 33793 2635
rect 32088 2604 33793 2632
rect 32088 2592 32094 2604
rect 33781 2601 33793 2604
rect 33827 2601 33839 2635
rect 33781 2595 33839 2601
rect 30558 2524 30564 2576
rect 30616 2564 30622 2576
rect 32309 2567 32367 2573
rect 32309 2564 32321 2567
rect 30616 2536 32321 2564
rect 30616 2524 30622 2536
rect 32309 2533 32321 2536
rect 32355 2533 32367 2567
rect 32309 2527 32367 2533
rect 33502 2524 33508 2576
rect 33560 2564 33566 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 33560 2536 34897 2564
rect 33560 2524 33566 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 34974 2524 34980 2576
rect 35032 2564 35038 2576
rect 36357 2567 36415 2573
rect 36357 2564 36369 2567
rect 35032 2536 36369 2564
rect 35032 2524 35038 2536
rect 36357 2533 36369 2536
rect 36403 2533 36415 2567
rect 36357 2527 36415 2533
rect 27249 2499 27307 2505
rect 27249 2465 27261 2499
rect 27295 2465 27307 2499
rect 30834 2496 30840 2508
rect 27249 2459 27307 2465
rect 28276 2468 30840 2496
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 22060 2400 22109 2428
rect 22060 2388 22066 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 22186 2388 22192 2440
rect 22244 2428 22250 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22244 2400 22385 2428
rect 22244 2388 22250 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 24854 2428 24860 2440
rect 23615 2400 24860 2428
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 24854 2388 24860 2400
rect 24912 2388 24918 2440
rect 24949 2431 25007 2437
rect 24949 2397 24961 2431
rect 24995 2397 25007 2431
rect 24949 2391 25007 2397
rect 19536 2360 19564 2388
rect 20349 2363 20407 2369
rect 20349 2360 20361 2363
rect 15120 2332 18644 2360
rect 19536 2332 20361 2360
rect 15930 2292 15936 2304
rect 14660 2264 15936 2292
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 16025 2295 16083 2301
rect 16025 2261 16037 2295
rect 16071 2292 16083 2295
rect 16482 2292 16488 2304
rect 16071 2264 16488 2292
rect 16071 2261 16083 2264
rect 16025 2255 16083 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 18616 2292 18644 2332
rect 20349 2329 20361 2332
rect 20395 2329 20407 2363
rect 24302 2360 24308 2372
rect 20349 2323 20407 2329
rect 20456 2332 24308 2360
rect 20456 2292 20484 2332
rect 24302 2320 24308 2332
rect 24360 2320 24366 2372
rect 24964 2360 24992 2391
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25556 2400 25605 2428
rect 25556 2388 25562 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 28276 2437 28304 2468
rect 30834 2456 30840 2468
rect 30892 2456 30898 2508
rect 34422 2496 34428 2508
rect 32140 2468 34428 2496
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28261 2431 28319 2437
rect 28261 2397 28273 2431
rect 28307 2397 28319 2431
rect 28261 2391 28319 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 28408 2400 29561 2428
rect 28408 2388 28414 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30374 2428 30380 2440
rect 30331 2400 30380 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 31018 2428 31024 2440
rect 30979 2400 31024 2428
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 32140 2437 32168 2468
rect 34422 2456 34428 2468
rect 34480 2456 34486 2508
rect 35986 2496 35992 2508
rect 34716 2468 35992 2496
rect 32125 2431 32183 2437
rect 32125 2397 32137 2431
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 32907 2400 33088 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 26234 2360 26240 2372
rect 24964 2332 26240 2360
rect 26234 2320 26240 2332
rect 26292 2320 26298 2372
rect 26878 2320 26884 2372
rect 26936 2360 26942 2372
rect 33060 2360 33088 2400
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 34716 2437 34744 2468
rect 35986 2456 35992 2468
rect 36044 2456 36050 2508
rect 37090 2496 37096 2508
rect 36096 2468 37096 2496
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33192 2400 33609 2428
rect 33192 2388 33198 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34701 2431 34759 2437
rect 34701 2397 34713 2431
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 35437 2431 35495 2437
rect 35437 2397 35449 2431
rect 35483 2428 35495 2431
rect 36096 2428 36124 2468
rect 37090 2456 37096 2468
rect 37148 2456 37154 2508
rect 35483 2400 36124 2428
rect 36173 2431 36231 2437
rect 35483 2397 35495 2400
rect 35437 2391 35495 2397
rect 36173 2397 36185 2431
rect 36219 2428 36231 2431
rect 36354 2428 36360 2440
rect 36219 2400 36360 2428
rect 36219 2397 36231 2400
rect 36173 2391 36231 2397
rect 36354 2388 36360 2400
rect 36412 2388 36418 2440
rect 35526 2360 35532 2372
rect 26936 2332 29776 2360
rect 33060 2332 35532 2360
rect 26936 2320 26942 2332
rect 18616 2264 20484 2292
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 21177 2295 21235 2301
rect 21177 2292 21189 2295
rect 20680 2264 21189 2292
rect 20680 2252 20686 2264
rect 21177 2261 21189 2264
rect 21223 2261 21235 2295
rect 21177 2255 21235 2261
rect 23753 2295 23811 2301
rect 23753 2261 23765 2295
rect 23799 2292 23811 2295
rect 23842 2292 23848 2304
rect 23799 2264 23848 2292
rect 23799 2261 23811 2264
rect 23753 2255 23811 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 26050 2252 26056 2304
rect 26108 2292 26114 2304
rect 29748 2301 29776 2332
rect 35526 2320 35532 2332
rect 35584 2320 35590 2372
rect 37921 2363 37979 2369
rect 37921 2329 37933 2363
rect 37967 2360 37979 2363
rect 39758 2360 39764 2372
rect 37967 2332 39764 2360
rect 37967 2329 37979 2332
rect 37921 2323 37979 2329
rect 39758 2320 39764 2332
rect 39816 2320 39822 2372
rect 28445 2295 28503 2301
rect 28445 2292 28457 2295
rect 26108 2264 28457 2292
rect 26108 2252 26114 2264
rect 28445 2261 28457 2264
rect 28491 2261 28503 2295
rect 28445 2255 28503 2261
rect 29733 2295 29791 2301
rect 29733 2261 29745 2295
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 29822 2252 29828 2304
rect 29880 2292 29886 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 29880 2264 31217 2292
rect 29880 2252 29886 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 33045 2295 33103 2301
rect 33045 2292 33057 2295
rect 31352 2264 33057 2292
rect 31352 2252 31358 2264
rect 33045 2261 33057 2264
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 34238 2252 34244 2304
rect 34296 2292 34302 2304
rect 35621 2295 35679 2301
rect 35621 2292 35633 2295
rect 34296 2264 35633 2292
rect 34296 2252 34302 2264
rect 35621 2261 35633 2264
rect 35667 2261 35679 2295
rect 38010 2292 38016 2304
rect 37971 2264 38016 2292
rect 35621 2255 35679 2261
rect 38010 2252 38016 2264
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 4614 2088 4620 2100
rect 3384 2060 4620 2088
rect 3384 2048 3390 2060
rect 4614 2048 4620 2060
rect 4672 2048 4678 2100
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 13262 2088 13268 2100
rect 5224 2060 13268 2088
rect 5224 2048 5230 2060
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 16390 2048 16396 2100
rect 16448 2088 16454 2100
rect 22186 2088 22192 2100
rect 16448 2060 22192 2088
rect 16448 2048 16454 2060
rect 22186 2048 22192 2060
rect 22244 2048 22250 2100
rect 30926 2088 30932 2100
rect 22388 2060 30932 2088
rect 2498 1980 2504 2032
rect 2556 2020 2562 2032
rect 9398 2020 9404 2032
rect 2556 1992 9404 2020
rect 2556 1980 2562 1992
rect 9398 1980 9404 1992
rect 9456 1980 9462 2032
rect 12250 1980 12256 2032
rect 12308 2020 12314 2032
rect 12308 1992 16344 2020
rect 12308 1980 12314 1992
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 3844 1924 12434 1952
rect 3844 1912 3850 1924
rect 3050 1844 3056 1896
rect 3108 1884 3114 1896
rect 10502 1884 10508 1896
rect 3108 1856 10508 1884
rect 3108 1844 3114 1856
rect 10502 1844 10508 1856
rect 10560 1844 10566 1896
rect 2406 1776 2412 1828
rect 2464 1816 2470 1828
rect 7190 1816 7196 1828
rect 2464 1788 7196 1816
rect 2464 1776 2470 1788
rect 7190 1776 7196 1788
rect 7248 1776 7254 1828
rect 12406 1816 12434 1924
rect 16316 1884 16344 1992
rect 18598 1980 18604 2032
rect 18656 2020 18662 2032
rect 22388 2020 22416 2060
rect 30926 2048 30932 2060
rect 30984 2048 30990 2100
rect 38010 2020 38016 2032
rect 18656 1992 22416 2020
rect 26206 1992 38016 2020
rect 18656 1980 18662 1992
rect 19794 1912 19800 1964
rect 19852 1952 19858 1964
rect 21266 1952 21272 1964
rect 19852 1924 21272 1952
rect 19852 1912 19858 1924
rect 21266 1912 21272 1924
rect 21324 1912 21330 1964
rect 21450 1912 21456 1964
rect 21508 1952 21514 1964
rect 26206 1952 26234 1992
rect 38010 1980 38016 1992
rect 38068 1980 38074 2032
rect 21508 1924 26234 1952
rect 21508 1912 21514 1924
rect 20438 1884 20444 1896
rect 16316 1856 20444 1884
rect 20438 1844 20444 1856
rect 20496 1844 20502 1896
rect 21358 1816 21364 1828
rect 12406 1788 21364 1816
rect 21358 1776 21364 1788
rect 21416 1776 21422 1828
rect 18322 1708 18328 1760
rect 18380 1748 18386 1760
rect 22094 1748 22100 1760
rect 18380 1720 22100 1748
rect 18380 1708 18386 1720
rect 22094 1708 22100 1720
rect 22152 1708 22158 1760
rect 3970 1504 3976 1556
rect 4028 1544 4034 1556
rect 5350 1544 5356 1556
rect 4028 1516 5356 1544
rect 4028 1504 4034 1516
rect 5350 1504 5356 1516
rect 5408 1504 5414 1556
rect 1854 1368 1860 1420
rect 1912 1408 1918 1420
rect 7926 1408 7932 1420
rect 1912 1380 7932 1408
rect 1912 1368 1918 1380
rect 7926 1368 7932 1380
rect 7984 1368 7990 1420
rect 17954 1368 17960 1420
rect 18012 1408 18018 1420
rect 20622 1408 20628 1420
rect 18012 1380 20628 1408
rect 18012 1368 18018 1380
rect 20622 1368 20628 1380
rect 20680 1368 20686 1420
rect 28350 1368 28356 1420
rect 28408 1408 28414 1420
rect 29822 1408 29828 1420
rect 28408 1380 29828 1408
rect 28408 1368 28414 1380
rect 29822 1368 29828 1380
rect 29880 1368 29886 1420
rect 2774 1232 2780 1284
rect 2832 1272 2838 1284
rect 4246 1272 4252 1284
rect 2832 1244 4252 1272
rect 2832 1232 2838 1244
rect 4246 1232 4252 1244
rect 4304 1232 4310 1284
rect 2590 1096 2596 1148
rect 2648 1136 2654 1148
rect 9030 1136 9036 1148
rect 2648 1108 9036 1136
rect 2648 1096 2654 1108
rect 9030 1096 9036 1108
rect 9088 1096 9094 1148
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 15200 47243 15252 47252
rect 15200 47209 15209 47243
rect 15209 47209 15243 47243
rect 15243 47209 15252 47243
rect 15200 47200 15252 47209
rect 25228 47243 25280 47252
rect 25228 47209 25237 47243
rect 25237 47209 25271 47243
rect 25271 47209 25280 47243
rect 25228 47200 25280 47209
rect 35348 47200 35400 47252
rect 5080 47039 5132 47048
rect 5080 47005 5089 47039
rect 5089 47005 5123 47039
rect 5123 47005 5132 47039
rect 5080 46996 5132 47005
rect 19248 46996 19300 47048
rect 24860 46996 24912 47048
rect 35348 46996 35400 47048
rect 5264 46903 5316 46912
rect 5264 46869 5273 46903
rect 5273 46869 5307 46903
rect 5307 46869 5316 46903
rect 5264 46860 5316 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 19248 46656 19300 46708
rect 20536 46520 20588 46572
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 20996 30676 21048 30728
rect 19248 30583 19300 30592
rect 19248 30549 19257 30583
rect 19257 30549 19291 30583
rect 19291 30549 19300 30583
rect 19248 30540 19300 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19248 30311 19300 30320
rect 15752 30200 15804 30252
rect 18420 30200 18472 30252
rect 19248 30277 19282 30311
rect 19282 30277 19300 30311
rect 19248 30268 19300 30277
rect 18512 30039 18564 30048
rect 18512 30005 18521 30039
rect 18521 30005 18555 30039
rect 18555 30005 18564 30039
rect 18512 29996 18564 30005
rect 20444 29996 20496 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 18420 29835 18472 29844
rect 18420 29801 18429 29835
rect 18429 29801 18463 29835
rect 18463 29801 18472 29835
rect 18420 29792 18472 29801
rect 20996 29835 21048 29844
rect 20996 29801 21005 29835
rect 21005 29801 21039 29835
rect 21039 29801 21048 29835
rect 20996 29792 21048 29801
rect 15752 29699 15804 29708
rect 15752 29665 15761 29699
rect 15761 29665 15795 29699
rect 15795 29665 15804 29699
rect 15752 29656 15804 29665
rect 20628 29699 20680 29708
rect 20628 29665 20637 29699
rect 20637 29665 20671 29699
rect 20671 29665 20680 29699
rect 20628 29656 20680 29665
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 17776 29631 17828 29640
rect 17776 29597 17785 29631
rect 17785 29597 17819 29631
rect 17819 29597 17828 29631
rect 17776 29588 17828 29597
rect 19984 29631 20036 29640
rect 19984 29597 19993 29631
rect 19993 29597 20027 29631
rect 20027 29597 20036 29631
rect 19984 29588 20036 29597
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 16672 29520 16724 29572
rect 17408 29452 17460 29504
rect 21272 29452 21324 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 16672 29291 16724 29300
rect 16672 29257 16681 29291
rect 16681 29257 16715 29291
rect 16715 29257 16724 29291
rect 16672 29248 16724 29257
rect 17776 29248 17828 29300
rect 20812 29248 20864 29300
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 18052 29155 18104 29164
rect 18052 29121 18061 29155
rect 18061 29121 18095 29155
rect 18095 29121 18104 29155
rect 18052 29112 18104 29121
rect 17960 29044 18012 29096
rect 19064 29155 19116 29164
rect 19064 29121 19073 29155
rect 19073 29121 19107 29155
rect 19107 29121 19116 29155
rect 19064 29112 19116 29121
rect 19248 29155 19300 29164
rect 18420 29044 18472 29096
rect 19248 29121 19257 29155
rect 19257 29121 19291 29155
rect 19291 29121 19300 29155
rect 19248 29112 19300 29121
rect 20444 29112 20496 29164
rect 22652 29112 22704 29164
rect 19892 29087 19944 29096
rect 19892 29053 19901 29087
rect 19901 29053 19935 29087
rect 19935 29053 19944 29087
rect 19892 29044 19944 29053
rect 18512 28976 18564 29028
rect 19156 28976 19208 29028
rect 16120 28908 16172 28960
rect 20812 28908 20864 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19984 28704 20036 28756
rect 20628 28704 20680 28756
rect 22652 28747 22704 28756
rect 15752 28568 15804 28620
rect 16120 28543 16172 28552
rect 16120 28509 16154 28543
rect 16154 28509 16172 28543
rect 16120 28500 16172 28509
rect 17960 28568 18012 28620
rect 22652 28713 22661 28747
rect 22661 28713 22695 28747
rect 22695 28713 22704 28747
rect 22652 28704 22704 28713
rect 18144 28500 18196 28552
rect 19340 28500 19392 28552
rect 19892 28500 19944 28552
rect 22100 28500 22152 28552
rect 17868 28475 17920 28484
rect 17868 28441 17877 28475
rect 17877 28441 17911 28475
rect 17911 28441 17920 28475
rect 17868 28432 17920 28441
rect 18788 28432 18840 28484
rect 19432 28475 19484 28484
rect 19432 28441 19441 28475
rect 19441 28441 19475 28475
rect 19475 28441 19484 28475
rect 19432 28432 19484 28441
rect 19984 28432 20036 28484
rect 21088 28432 21140 28484
rect 18236 28407 18288 28416
rect 18236 28373 18245 28407
rect 18245 28373 18279 28407
rect 18279 28373 18288 28407
rect 18236 28364 18288 28373
rect 20628 28364 20680 28416
rect 21824 28407 21876 28416
rect 21824 28373 21833 28407
rect 21833 28373 21867 28407
rect 21867 28373 21876 28407
rect 21824 28364 21876 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 15936 28160 15988 28212
rect 16856 28160 16908 28212
rect 17868 28160 17920 28212
rect 18052 28160 18104 28212
rect 19248 28160 19300 28212
rect 20628 28203 20680 28212
rect 20628 28169 20637 28203
rect 20637 28169 20671 28203
rect 20671 28169 20680 28203
rect 20628 28160 20680 28169
rect 21088 28203 21140 28212
rect 21088 28169 21097 28203
rect 21097 28169 21131 28203
rect 21131 28169 21140 28203
rect 21088 28160 21140 28169
rect 15384 28024 15436 28076
rect 18236 28092 18288 28144
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 15292 27956 15344 28008
rect 17592 27956 17644 28008
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 19156 27956 19208 28008
rect 17960 27888 18012 27940
rect 20260 28067 20312 28076
rect 20260 28033 20269 28067
rect 20269 28033 20303 28067
rect 20303 28033 20312 28067
rect 20260 28024 20312 28033
rect 21272 28067 21324 28076
rect 20168 27956 20220 28008
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 21364 28024 21416 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 22100 28024 22152 28076
rect 24400 28024 24452 28076
rect 20812 27956 20864 28008
rect 25136 28024 25188 28076
rect 18788 27820 18840 27872
rect 21824 27863 21876 27872
rect 21824 27829 21833 27863
rect 21833 27829 21867 27863
rect 21867 27829 21876 27863
rect 21824 27820 21876 27829
rect 24216 27820 24268 27872
rect 24768 27820 24820 27872
rect 26056 27820 26108 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 20260 27616 20312 27668
rect 18144 27548 18196 27600
rect 19432 27548 19484 27600
rect 24400 27591 24452 27600
rect 24400 27557 24409 27591
rect 24409 27557 24443 27591
rect 24443 27557 24452 27591
rect 24400 27548 24452 27557
rect 15476 27480 15528 27532
rect 17040 27480 17092 27532
rect 19340 27480 19392 27532
rect 21824 27480 21876 27532
rect 22100 27523 22152 27532
rect 22100 27489 22109 27523
rect 22109 27489 22143 27523
rect 22143 27489 22152 27523
rect 22100 27480 22152 27489
rect 15752 27412 15804 27464
rect 13360 27344 13412 27396
rect 12440 27276 12492 27328
rect 15292 27344 15344 27396
rect 17500 27412 17552 27464
rect 18052 27412 18104 27464
rect 19156 27412 19208 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 25228 27455 25280 27464
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 22376 27387 22428 27396
rect 22376 27353 22410 27387
rect 22410 27353 22428 27387
rect 22376 27344 22428 27353
rect 14924 27276 14976 27328
rect 19984 27276 20036 27328
rect 20812 27319 20864 27328
rect 20812 27285 20821 27319
rect 20821 27285 20855 27319
rect 20855 27285 20864 27319
rect 20812 27276 20864 27285
rect 21272 27276 21324 27328
rect 22560 27276 22612 27328
rect 25320 27319 25372 27328
rect 25320 27285 25329 27319
rect 25329 27285 25363 27319
rect 25363 27285 25372 27319
rect 25320 27276 25372 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 13360 27115 13412 27124
rect 13360 27081 13369 27115
rect 13369 27081 13403 27115
rect 13403 27081 13412 27115
rect 13360 27072 13412 27081
rect 16856 27072 16908 27124
rect 19064 27072 19116 27124
rect 20168 27072 20220 27124
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 15752 27004 15804 27056
rect 17408 27004 17460 27056
rect 17960 27004 18012 27056
rect 16212 26936 16264 26988
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 19156 27004 19208 27056
rect 19800 27004 19852 27056
rect 20260 26936 20312 26988
rect 20720 26936 20772 26988
rect 25228 27004 25280 27056
rect 22560 26979 22612 26988
rect 21640 26868 21692 26920
rect 22560 26945 22569 26979
rect 22569 26945 22603 26979
rect 22603 26945 22612 26979
rect 22560 26936 22612 26945
rect 26240 27004 26292 27056
rect 20352 26800 20404 26852
rect 21824 26800 21876 26852
rect 26056 26979 26108 26988
rect 23848 26868 23900 26920
rect 24216 26911 24268 26920
rect 24216 26877 24225 26911
rect 24225 26877 24259 26911
rect 24259 26877 24268 26911
rect 24216 26868 24268 26877
rect 24768 26868 24820 26920
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 26884 26936 26936 26988
rect 24032 26843 24084 26852
rect 15936 26732 15988 26784
rect 16028 26775 16080 26784
rect 16028 26741 16037 26775
rect 16037 26741 16071 26775
rect 16071 26741 16080 26775
rect 23756 26775 23808 26784
rect 16028 26732 16080 26741
rect 23756 26741 23765 26775
rect 23765 26741 23799 26775
rect 23799 26741 23808 26775
rect 23756 26732 23808 26741
rect 24032 26809 24041 26843
rect 24041 26809 24075 26843
rect 24075 26809 24084 26843
rect 24032 26800 24084 26809
rect 25228 26800 25280 26852
rect 26424 26800 26476 26852
rect 25044 26732 25096 26784
rect 25596 26732 25648 26784
rect 27620 26732 27672 26784
rect 27896 26732 27948 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 14188 26528 14240 26580
rect 15936 26528 15988 26580
rect 16856 26528 16908 26580
rect 18328 26528 18380 26580
rect 19340 26571 19392 26580
rect 19340 26537 19349 26571
rect 19349 26537 19383 26571
rect 19383 26537 19392 26571
rect 19340 26528 19392 26537
rect 20904 26528 20956 26580
rect 22192 26571 22244 26580
rect 22192 26537 22201 26571
rect 22201 26537 22235 26571
rect 22235 26537 22244 26571
rect 22192 26528 22244 26537
rect 23848 26571 23900 26580
rect 19248 26460 19300 26512
rect 12440 26324 12492 26376
rect 13636 26324 13688 26376
rect 13084 26256 13136 26308
rect 15016 26324 15068 26376
rect 14464 26299 14516 26308
rect 14464 26265 14473 26299
rect 14473 26265 14507 26299
rect 14507 26265 14516 26299
rect 14464 26256 14516 26265
rect 14924 26256 14976 26308
rect 15936 26324 15988 26376
rect 19064 26392 19116 26444
rect 15660 26256 15712 26308
rect 18236 26324 18288 26376
rect 19340 26367 19392 26376
rect 17408 26299 17460 26308
rect 17408 26265 17417 26299
rect 17417 26265 17451 26299
rect 17451 26265 17460 26299
rect 17408 26256 17460 26265
rect 17500 26299 17552 26308
rect 17500 26265 17509 26299
rect 17509 26265 17543 26299
rect 17543 26265 17552 26299
rect 17500 26256 17552 26265
rect 18604 26256 18656 26308
rect 19340 26333 19349 26367
rect 19349 26333 19383 26367
rect 19383 26333 19392 26367
rect 19340 26324 19392 26333
rect 19800 26324 19852 26376
rect 22652 26460 22704 26512
rect 23848 26537 23857 26571
rect 23857 26537 23891 26571
rect 23891 26537 23900 26571
rect 23848 26528 23900 26537
rect 24032 26528 24084 26580
rect 25136 26571 25188 26580
rect 25136 26537 25145 26571
rect 25145 26537 25179 26571
rect 25179 26537 25188 26571
rect 25136 26528 25188 26537
rect 26884 26571 26936 26580
rect 26884 26537 26893 26571
rect 26893 26537 26927 26571
rect 26927 26537 26936 26571
rect 26884 26528 26936 26537
rect 24216 26460 24268 26512
rect 25228 26460 25280 26512
rect 20168 26324 20220 26376
rect 20444 26324 20496 26376
rect 21640 26324 21692 26376
rect 22560 26324 22612 26376
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 25780 26367 25832 26376
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 26240 26367 26292 26376
rect 25780 26324 25832 26333
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26424 26367 26476 26376
rect 26424 26333 26433 26367
rect 26433 26333 26467 26367
rect 26467 26333 26476 26367
rect 26424 26324 26476 26333
rect 27068 26367 27120 26376
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 13176 26231 13228 26240
rect 13176 26197 13185 26231
rect 13185 26197 13219 26231
rect 13219 26197 13228 26231
rect 13176 26188 13228 26197
rect 15292 26188 15344 26240
rect 23112 26256 23164 26308
rect 23572 26256 23624 26308
rect 26516 26256 26568 26308
rect 27712 26324 27764 26376
rect 27896 26367 27948 26376
rect 27896 26333 27906 26367
rect 27906 26333 27940 26367
rect 27940 26333 27948 26367
rect 27896 26324 27948 26333
rect 27988 26367 28040 26376
rect 27988 26333 27997 26367
rect 27997 26333 28031 26367
rect 28031 26333 28040 26367
rect 27988 26324 28040 26333
rect 27804 26256 27856 26308
rect 22008 26188 22060 26240
rect 22652 26188 22704 26240
rect 28080 26188 28132 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 14464 25984 14516 26036
rect 14740 25916 14792 25968
rect 15936 25916 15988 25968
rect 18696 25916 18748 25968
rect 12256 25848 12308 25900
rect 14924 25848 14976 25900
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 18604 25891 18656 25900
rect 11796 25780 11848 25832
rect 15476 25780 15528 25832
rect 15660 25780 15712 25832
rect 18604 25857 18613 25891
rect 18613 25857 18647 25891
rect 18647 25857 18656 25891
rect 18604 25848 18656 25857
rect 20076 25984 20128 26036
rect 21364 25984 21416 26036
rect 25320 25984 25372 26036
rect 20076 25891 20128 25900
rect 18512 25780 18564 25832
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 20812 25891 20864 25900
rect 20812 25857 20821 25891
rect 20821 25857 20855 25891
rect 20855 25857 20864 25891
rect 20812 25848 20864 25857
rect 22744 25916 22796 25968
rect 27068 25984 27120 26036
rect 20720 25780 20772 25832
rect 21272 25780 21324 25832
rect 22560 25848 22612 25900
rect 22836 25891 22888 25900
rect 22836 25857 22845 25891
rect 22845 25857 22879 25891
rect 22879 25857 22888 25891
rect 22836 25848 22888 25857
rect 24308 25891 24360 25900
rect 24308 25857 24317 25891
rect 24317 25857 24351 25891
rect 24351 25857 24360 25891
rect 24308 25848 24360 25857
rect 25320 25891 25372 25900
rect 23112 25780 23164 25832
rect 25320 25857 25329 25891
rect 25329 25857 25363 25891
rect 25363 25857 25372 25891
rect 25320 25848 25372 25857
rect 26240 25891 26292 25900
rect 24768 25780 24820 25832
rect 25412 25712 25464 25764
rect 26240 25857 26249 25891
rect 26249 25857 26283 25891
rect 26283 25857 26292 25891
rect 26240 25848 26292 25857
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 28632 25916 28684 25968
rect 27896 25848 27948 25900
rect 28080 25891 28132 25900
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 28264 25848 28316 25900
rect 26792 25780 26844 25832
rect 27712 25780 27764 25832
rect 30564 25848 30616 25900
rect 29368 25780 29420 25832
rect 34796 25780 34848 25832
rect 27804 25755 27856 25764
rect 27804 25721 27813 25755
rect 27813 25721 27847 25755
rect 27847 25721 27856 25755
rect 27804 25712 27856 25721
rect 13268 25644 13320 25696
rect 17500 25687 17552 25696
rect 17500 25653 17509 25687
rect 17509 25653 17543 25687
rect 17543 25653 17552 25687
rect 17500 25644 17552 25653
rect 18420 25687 18472 25696
rect 18420 25653 18429 25687
rect 18429 25653 18463 25687
rect 18463 25653 18472 25687
rect 18420 25644 18472 25653
rect 19892 25687 19944 25696
rect 19892 25653 19901 25687
rect 19901 25653 19935 25687
rect 19935 25653 19944 25687
rect 19892 25644 19944 25653
rect 20904 25644 20956 25696
rect 22468 25644 22520 25696
rect 25688 25644 25740 25696
rect 27896 25644 27948 25696
rect 32864 25644 32916 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 12256 25440 12308 25492
rect 5264 25304 5316 25356
rect 19892 25440 19944 25492
rect 20904 25440 20956 25492
rect 24584 25440 24636 25492
rect 24768 25440 24820 25492
rect 18052 25372 18104 25424
rect 20720 25415 20772 25424
rect 20720 25381 20729 25415
rect 20729 25381 20763 25415
rect 20763 25381 20772 25415
rect 20720 25372 20772 25381
rect 13176 25236 13228 25288
rect 15292 25304 15344 25356
rect 15752 25304 15804 25356
rect 16304 25347 16356 25356
rect 16304 25313 16313 25347
rect 16313 25313 16347 25347
rect 16347 25313 16356 25347
rect 16304 25304 16356 25313
rect 14740 25236 14792 25288
rect 17500 25236 17552 25288
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 20260 25304 20312 25356
rect 21272 25372 21324 25424
rect 22468 25304 22520 25356
rect 22560 25347 22612 25356
rect 22560 25313 22569 25347
rect 22569 25313 22603 25347
rect 22603 25313 22612 25347
rect 23020 25347 23072 25356
rect 22560 25304 22612 25313
rect 23020 25313 23029 25347
rect 23029 25313 23063 25347
rect 23063 25313 23072 25347
rect 23020 25304 23072 25313
rect 24860 25304 24912 25356
rect 19432 25279 19484 25288
rect 19432 25245 19435 25279
rect 19435 25245 19469 25279
rect 19469 25245 19484 25279
rect 19432 25236 19484 25245
rect 20812 25236 20864 25288
rect 23112 25236 23164 25288
rect 23756 25236 23808 25288
rect 25136 25279 25188 25288
rect 20720 25168 20772 25220
rect 23940 25168 23992 25220
rect 25136 25245 25145 25279
rect 25145 25245 25179 25279
rect 25179 25245 25188 25279
rect 25136 25236 25188 25245
rect 25688 25236 25740 25288
rect 27620 25279 27672 25288
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 27896 25279 27948 25288
rect 27896 25245 27930 25279
rect 27930 25245 27948 25279
rect 27896 25236 27948 25245
rect 29828 25279 29880 25288
rect 29828 25245 29837 25279
rect 29837 25245 29871 25279
rect 29871 25245 29880 25279
rect 31668 25279 31720 25288
rect 29828 25236 29880 25245
rect 31668 25245 31677 25279
rect 31677 25245 31711 25279
rect 31711 25245 31720 25279
rect 31668 25236 31720 25245
rect 25044 25168 25096 25220
rect 27160 25168 27212 25220
rect 30472 25168 30524 25220
rect 30748 25168 30800 25220
rect 12808 25143 12860 25152
rect 12808 25109 12817 25143
rect 12817 25109 12851 25143
rect 12851 25109 12860 25143
rect 12808 25100 12860 25109
rect 13176 25143 13228 25152
rect 13176 25109 13185 25143
rect 13185 25109 13219 25143
rect 13219 25109 13228 25143
rect 13176 25100 13228 25109
rect 17224 25100 17276 25152
rect 17960 25100 18012 25152
rect 26240 25100 26292 25152
rect 28172 25100 28224 25152
rect 31208 25143 31260 25152
rect 31208 25109 31217 25143
rect 31217 25109 31251 25143
rect 31251 25109 31260 25143
rect 31208 25100 31260 25109
rect 31300 25100 31352 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 17224 24896 17276 24948
rect 18696 24939 18748 24948
rect 18696 24905 18705 24939
rect 18705 24905 18739 24939
rect 18739 24905 18748 24939
rect 18696 24896 18748 24905
rect 12808 24828 12860 24880
rect 15200 24828 15252 24880
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 17868 24828 17920 24880
rect 23756 24896 23808 24948
rect 25136 24896 25188 24948
rect 13268 24692 13320 24744
rect 13360 24556 13412 24608
rect 14648 24692 14700 24744
rect 18052 24760 18104 24812
rect 15292 24735 15344 24744
rect 15292 24701 15301 24735
rect 15301 24701 15335 24735
rect 15335 24701 15344 24735
rect 15292 24692 15344 24701
rect 17132 24692 17184 24744
rect 17960 24692 18012 24744
rect 13636 24667 13688 24676
rect 13636 24633 13645 24667
rect 13645 24633 13679 24667
rect 13679 24633 13688 24667
rect 13636 24624 13688 24633
rect 18512 24803 18564 24812
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 19984 24760 20036 24812
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 20812 24803 20864 24812
rect 20812 24769 20821 24803
rect 20821 24769 20855 24803
rect 20855 24769 20864 24803
rect 20812 24760 20864 24769
rect 21548 24760 21600 24812
rect 23020 24760 23072 24812
rect 24216 24803 24268 24812
rect 24216 24769 24225 24803
rect 24225 24769 24259 24803
rect 24259 24769 24268 24803
rect 24216 24760 24268 24769
rect 24308 24760 24360 24812
rect 24768 24760 24820 24812
rect 26240 24939 26292 24948
rect 26240 24905 26265 24939
rect 26265 24905 26292 24939
rect 26240 24896 26292 24905
rect 27620 24896 27672 24948
rect 26148 24828 26200 24880
rect 18880 24692 18932 24744
rect 19248 24692 19300 24744
rect 21916 24692 21968 24744
rect 22468 24692 22520 24744
rect 26240 24760 26292 24812
rect 26792 24760 26844 24812
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 25596 24692 25648 24744
rect 15016 24556 15068 24608
rect 17500 24556 17552 24608
rect 18236 24556 18288 24608
rect 20628 24599 20680 24608
rect 20628 24565 20637 24599
rect 20637 24565 20671 24599
rect 20671 24565 20680 24599
rect 20628 24556 20680 24565
rect 20904 24624 20956 24676
rect 22836 24624 22888 24676
rect 25228 24667 25280 24676
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 24032 24599 24084 24608
rect 24032 24565 24041 24599
rect 24041 24565 24075 24599
rect 24075 24565 24084 24599
rect 24032 24556 24084 24565
rect 25228 24633 25237 24667
rect 25237 24633 25271 24667
rect 25271 24633 25280 24667
rect 25228 24624 25280 24633
rect 26332 24624 26384 24676
rect 27712 24760 27764 24812
rect 27988 24760 28040 24812
rect 27896 24624 27948 24676
rect 26516 24556 26568 24608
rect 27068 24599 27120 24608
rect 27068 24565 27077 24599
rect 27077 24565 27111 24599
rect 27111 24565 27120 24599
rect 27068 24556 27120 24565
rect 27712 24556 27764 24608
rect 28540 24803 28592 24812
rect 28540 24769 28549 24803
rect 28549 24769 28583 24803
rect 28583 24769 28592 24803
rect 29828 24828 29880 24880
rect 28540 24760 28592 24769
rect 30380 24760 30432 24812
rect 32680 24760 32732 24812
rect 29000 24556 29052 24608
rect 29828 24556 29880 24608
rect 32036 24692 32088 24744
rect 30288 24624 30340 24676
rect 32312 24556 32364 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 16856 24352 16908 24404
rect 20628 24352 20680 24404
rect 21824 24352 21876 24404
rect 24216 24352 24268 24404
rect 26240 24352 26292 24404
rect 27804 24352 27856 24404
rect 15200 24284 15252 24336
rect 16028 24284 16080 24336
rect 15016 24259 15068 24268
rect 15016 24225 15025 24259
rect 15025 24225 15059 24259
rect 15059 24225 15068 24259
rect 15016 24216 15068 24225
rect 18328 24284 18380 24336
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 13084 24148 13136 24200
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 13176 24123 13228 24132
rect 13176 24089 13185 24123
rect 13185 24089 13219 24123
rect 13219 24089 13228 24123
rect 13176 24080 13228 24089
rect 13452 24080 13504 24132
rect 16488 24148 16540 24200
rect 16948 24148 17000 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 18880 24216 18932 24268
rect 16580 24080 16632 24132
rect 17040 24080 17092 24132
rect 17224 24080 17276 24132
rect 17776 24148 17828 24200
rect 19340 24216 19392 24268
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 19892 24191 19944 24200
rect 19892 24157 19901 24191
rect 19901 24157 19935 24191
rect 19935 24157 19944 24191
rect 19892 24148 19944 24157
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 21548 24216 21600 24268
rect 22192 24216 22244 24268
rect 22468 24216 22520 24268
rect 24124 24216 24176 24268
rect 32772 24352 32824 24404
rect 34704 24352 34756 24404
rect 31208 24216 31260 24268
rect 20812 24148 20864 24200
rect 22008 24191 22060 24200
rect 22008 24157 22017 24191
rect 22017 24157 22051 24191
rect 22051 24157 22060 24191
rect 22008 24148 22060 24157
rect 24032 24148 24084 24200
rect 19156 24080 19208 24132
rect 24676 24148 24728 24200
rect 27436 24191 27488 24200
rect 26056 24080 26108 24132
rect 27436 24157 27445 24191
rect 27445 24157 27479 24191
rect 27479 24157 27488 24191
rect 27436 24148 27488 24157
rect 27712 24191 27764 24200
rect 27712 24157 27746 24191
rect 27746 24157 27764 24191
rect 27712 24148 27764 24157
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 30932 24191 30984 24200
rect 28448 24080 28500 24132
rect 30932 24157 30941 24191
rect 30941 24157 30975 24191
rect 30975 24157 30984 24191
rect 30932 24148 30984 24157
rect 31668 24148 31720 24200
rect 30840 24080 30892 24132
rect 31300 24080 31352 24132
rect 32956 24080 33008 24132
rect 33048 24080 33100 24132
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 12900 24012 12952 24064
rect 18236 24012 18288 24064
rect 18512 24012 18564 24064
rect 19984 24055 20036 24064
rect 19984 24021 19993 24055
rect 19993 24021 20027 24055
rect 20027 24021 20036 24055
rect 19984 24012 20036 24021
rect 20168 24012 20220 24064
rect 25596 24055 25648 24064
rect 25596 24021 25621 24055
rect 25621 24021 25648 24055
rect 25780 24055 25832 24064
rect 25596 24012 25648 24021
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 27712 24012 27764 24064
rect 27896 24012 27948 24064
rect 28356 24012 28408 24064
rect 28540 24012 28592 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 13176 23808 13228 23860
rect 12348 23740 12400 23792
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 13452 23536 13504 23588
rect 15844 23808 15896 23860
rect 16764 23808 16816 23860
rect 18604 23808 18656 23860
rect 21916 23808 21968 23860
rect 24308 23808 24360 23860
rect 24768 23808 24820 23860
rect 19984 23740 20036 23792
rect 20076 23740 20128 23792
rect 15660 23672 15712 23724
rect 16212 23672 16264 23724
rect 17868 23715 17920 23724
rect 15568 23647 15620 23656
rect 15568 23613 15577 23647
rect 15577 23613 15611 23647
rect 15611 23613 15620 23647
rect 15568 23604 15620 23613
rect 16948 23604 17000 23656
rect 17868 23681 17877 23715
rect 17877 23681 17911 23715
rect 17911 23681 17920 23715
rect 17868 23672 17920 23681
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 18512 23672 18564 23724
rect 20168 23672 20220 23724
rect 14648 23536 14700 23588
rect 18420 23604 18472 23656
rect 19984 23604 20036 23656
rect 20444 23662 20496 23714
rect 20720 23672 20772 23724
rect 21272 23672 21324 23724
rect 21732 23672 21784 23724
rect 22192 23672 22244 23724
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 25320 23740 25372 23792
rect 25688 23740 25740 23792
rect 22836 23672 22888 23681
rect 21916 23604 21968 23656
rect 25504 23672 25556 23724
rect 25964 23715 26016 23724
rect 25964 23681 25973 23715
rect 25973 23681 26007 23715
rect 26007 23681 26016 23715
rect 25964 23672 26016 23681
rect 27988 23808 28040 23860
rect 28632 23808 28684 23860
rect 20444 23536 20496 23588
rect 23848 23579 23900 23588
rect 23848 23545 23857 23579
rect 23857 23545 23891 23579
rect 23891 23545 23900 23579
rect 23848 23536 23900 23545
rect 25044 23604 25096 23656
rect 29000 23783 29052 23792
rect 29000 23749 29009 23783
rect 29009 23749 29043 23783
rect 29043 23749 29052 23783
rect 29000 23740 29052 23749
rect 29920 23740 29972 23792
rect 30564 23740 30616 23792
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 16948 23468 17000 23520
rect 19524 23511 19576 23520
rect 19524 23477 19533 23511
rect 19533 23477 19567 23511
rect 19567 23477 19576 23511
rect 19524 23468 19576 23477
rect 20996 23468 21048 23520
rect 21824 23468 21876 23520
rect 22560 23468 22612 23520
rect 24308 23468 24360 23520
rect 24768 23468 24820 23520
rect 25228 23536 25280 23588
rect 28172 23672 28224 23724
rect 28356 23604 28408 23656
rect 28540 23647 28592 23656
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 29276 23715 29328 23724
rect 29276 23681 29285 23715
rect 29285 23681 29319 23715
rect 29319 23681 29328 23715
rect 29276 23672 29328 23681
rect 28540 23604 28592 23613
rect 28816 23536 28868 23588
rect 31760 23672 31812 23724
rect 30564 23647 30616 23656
rect 30564 23613 30573 23647
rect 30573 23613 30607 23647
rect 30607 23613 30616 23647
rect 30564 23604 30616 23613
rect 32956 23808 33008 23860
rect 33416 23808 33468 23860
rect 32036 23740 32088 23792
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32496 23740 32548 23792
rect 32772 23672 32824 23724
rect 32956 23672 33008 23724
rect 33784 23715 33836 23724
rect 33784 23681 33793 23715
rect 33793 23681 33827 23715
rect 33827 23681 33836 23715
rect 33784 23672 33836 23681
rect 34428 23715 34480 23724
rect 34428 23681 34437 23715
rect 34437 23681 34471 23715
rect 34471 23681 34480 23715
rect 34428 23672 34480 23681
rect 32772 23536 32824 23588
rect 32864 23536 32916 23588
rect 33784 23536 33836 23588
rect 34152 23604 34204 23656
rect 34428 23536 34480 23588
rect 28264 23468 28316 23520
rect 31392 23468 31444 23520
rect 32128 23468 32180 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 12440 23128 12492 23180
rect 16672 23264 16724 23316
rect 18052 23264 18104 23316
rect 12900 23060 12952 23112
rect 13084 23060 13136 23112
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 15660 23196 15712 23248
rect 16580 23196 16632 23248
rect 19616 23264 19668 23316
rect 20444 23307 20496 23316
rect 20444 23273 20453 23307
rect 20453 23273 20487 23307
rect 20487 23273 20496 23307
rect 20444 23264 20496 23273
rect 22928 23307 22980 23316
rect 22928 23273 22937 23307
rect 22937 23273 22971 23307
rect 22971 23273 22980 23307
rect 22928 23264 22980 23273
rect 26148 23264 26200 23316
rect 30472 23264 30524 23316
rect 34796 23307 34848 23316
rect 34796 23273 34805 23307
rect 34805 23273 34839 23307
rect 34839 23273 34848 23307
rect 34796 23264 34848 23273
rect 14832 23128 14884 23180
rect 16212 23128 16264 23180
rect 17040 23128 17092 23180
rect 18052 23128 18104 23180
rect 18328 23171 18380 23180
rect 18328 23137 18337 23171
rect 18337 23137 18371 23171
rect 18371 23137 18380 23171
rect 18328 23128 18380 23137
rect 13452 22992 13504 23044
rect 13084 22924 13136 22976
rect 13176 22924 13228 22976
rect 17592 23060 17644 23112
rect 18144 23060 18196 23112
rect 27068 23196 27120 23248
rect 27528 23239 27580 23248
rect 27528 23205 27537 23239
rect 27537 23205 27571 23239
rect 27571 23205 27580 23239
rect 27528 23196 27580 23205
rect 30380 23196 30432 23248
rect 19432 23128 19484 23180
rect 20168 23128 20220 23180
rect 20720 23128 20772 23180
rect 21180 23128 21232 23180
rect 19340 23060 19392 23112
rect 18604 22992 18656 23044
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 19892 23060 19944 23112
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 21824 23060 21876 23112
rect 23756 23128 23808 23180
rect 24032 23128 24084 23180
rect 24768 23128 24820 23180
rect 23204 23060 23256 23112
rect 16764 22924 16816 22976
rect 17316 22924 17368 22976
rect 17592 22924 17644 22976
rect 18328 22924 18380 22976
rect 22376 22924 22428 22976
rect 23572 22924 23624 22976
rect 23756 22992 23808 23044
rect 24860 23060 24912 23112
rect 29736 23128 29788 23180
rect 25596 23060 25648 23112
rect 30012 23060 30064 23112
rect 31024 23128 31076 23180
rect 32496 23171 32548 23180
rect 32496 23137 32505 23171
rect 32505 23137 32539 23171
rect 32539 23137 32548 23171
rect 32496 23128 32548 23137
rect 27160 23035 27212 23044
rect 23848 22924 23900 22976
rect 26056 22924 26108 22976
rect 27160 23001 27169 23035
rect 27169 23001 27203 23035
rect 27203 23001 27212 23035
rect 27160 22992 27212 23001
rect 27528 22992 27580 23044
rect 28632 23035 28684 23044
rect 28632 23001 28641 23035
rect 28641 23001 28675 23035
rect 28675 23001 28684 23035
rect 28632 22992 28684 23001
rect 30472 23103 30524 23112
rect 30472 23069 30481 23103
rect 30481 23069 30515 23103
rect 30515 23069 30524 23103
rect 30472 23060 30524 23069
rect 30932 23060 30984 23112
rect 31392 23103 31444 23112
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 32128 23103 32180 23112
rect 30380 22992 30432 23044
rect 30564 22992 30616 23044
rect 31208 22992 31260 23044
rect 32128 23069 32137 23103
rect 32137 23069 32171 23103
rect 32171 23069 32180 23103
rect 32128 23060 32180 23069
rect 32312 23103 32364 23112
rect 32312 23069 32321 23103
rect 32321 23069 32355 23103
rect 32355 23069 32364 23103
rect 32312 23060 32364 23069
rect 32404 23103 32456 23112
rect 32404 23069 32413 23103
rect 32413 23069 32447 23103
rect 32447 23069 32456 23103
rect 32956 23128 33008 23180
rect 32404 23060 32456 23069
rect 33324 23103 33376 23112
rect 33324 23069 33333 23103
rect 33333 23069 33367 23103
rect 33367 23069 33376 23103
rect 33324 23060 33376 23069
rect 34704 23103 34756 23112
rect 34704 23069 34713 23103
rect 34713 23069 34747 23103
rect 34747 23069 34756 23103
rect 34704 23060 34756 23069
rect 29644 22924 29696 22976
rect 30104 22924 30156 22976
rect 32864 22967 32916 22976
rect 32864 22933 32873 22967
rect 32873 22933 32907 22967
rect 32907 22933 32916 22967
rect 32864 22924 32916 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 14832 22763 14884 22772
rect 14832 22729 14841 22763
rect 14841 22729 14875 22763
rect 14875 22729 14884 22763
rect 14832 22720 14884 22729
rect 11796 22584 11848 22636
rect 12808 22652 12860 22704
rect 13084 22652 13136 22704
rect 14280 22516 14332 22568
rect 18328 22720 18380 22772
rect 15660 22652 15712 22704
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 16304 22584 16356 22636
rect 18236 22652 18288 22704
rect 19248 22652 19300 22704
rect 19340 22627 19392 22636
rect 19340 22593 19349 22627
rect 19349 22593 19383 22627
rect 19383 22593 19392 22627
rect 19340 22584 19392 22593
rect 17132 22516 17184 22568
rect 13452 22380 13504 22432
rect 16672 22448 16724 22500
rect 14464 22423 14516 22432
rect 14464 22389 14473 22423
rect 14473 22389 14507 22423
rect 14507 22389 14516 22423
rect 14464 22380 14516 22389
rect 15200 22380 15252 22432
rect 18604 22423 18656 22432
rect 18604 22389 18613 22423
rect 18613 22389 18647 22423
rect 18647 22389 18656 22423
rect 18604 22380 18656 22389
rect 21088 22720 21140 22772
rect 21272 22720 21324 22772
rect 20076 22584 20128 22636
rect 20628 22652 20680 22704
rect 22100 22652 22152 22704
rect 20904 22584 20956 22636
rect 20996 22584 21048 22636
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 21824 22584 21876 22636
rect 22376 22695 22428 22704
rect 22376 22661 22385 22695
rect 22385 22661 22419 22695
rect 22419 22661 22428 22695
rect 27344 22720 27396 22772
rect 28816 22763 28868 22772
rect 28816 22729 28825 22763
rect 28825 22729 28859 22763
rect 28859 22729 28868 22763
rect 28816 22720 28868 22729
rect 29736 22763 29788 22772
rect 29736 22729 29745 22763
rect 29745 22729 29779 22763
rect 29779 22729 29788 22763
rect 29736 22720 29788 22729
rect 29828 22720 29880 22772
rect 30564 22720 30616 22772
rect 30748 22720 30800 22772
rect 32404 22720 32456 22772
rect 22376 22652 22428 22661
rect 20260 22448 20312 22500
rect 19524 22380 19576 22432
rect 23848 22448 23900 22500
rect 25872 22652 25924 22704
rect 27528 22695 27580 22704
rect 27528 22661 27537 22695
rect 27537 22661 27571 22695
rect 27571 22661 27580 22695
rect 30104 22695 30156 22704
rect 27528 22652 27580 22661
rect 24952 22627 25004 22636
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 26148 22584 26200 22636
rect 27804 22584 27856 22636
rect 25504 22516 25556 22568
rect 26056 22516 26108 22568
rect 28080 22584 28132 22636
rect 28448 22584 28500 22636
rect 30104 22661 30113 22695
rect 30113 22661 30147 22695
rect 30147 22661 30156 22695
rect 30104 22652 30156 22661
rect 32036 22652 32088 22704
rect 32772 22652 32824 22704
rect 32864 22652 32916 22704
rect 29920 22627 29972 22636
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30840 22584 30892 22636
rect 31021 22627 31073 22636
rect 31021 22593 31030 22627
rect 31030 22593 31064 22627
rect 31064 22593 31073 22627
rect 31021 22584 31073 22593
rect 31116 22627 31168 22636
rect 31116 22593 31125 22627
rect 31125 22593 31159 22627
rect 31159 22593 31168 22627
rect 31116 22584 31168 22593
rect 30288 22516 30340 22568
rect 30748 22516 30800 22568
rect 31760 22584 31812 22636
rect 32312 22584 32364 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33140 22584 33192 22636
rect 33416 22584 33468 22636
rect 33232 22516 33284 22568
rect 25688 22448 25740 22500
rect 27804 22491 27856 22500
rect 27804 22457 27813 22491
rect 27813 22457 27847 22491
rect 27847 22457 27856 22491
rect 27804 22448 27856 22457
rect 27896 22491 27948 22500
rect 27896 22457 27905 22491
rect 27905 22457 27939 22491
rect 27939 22457 27948 22491
rect 27896 22448 27948 22457
rect 20720 22380 20772 22432
rect 22560 22423 22612 22432
rect 22560 22389 22569 22423
rect 22569 22389 22603 22423
rect 22603 22389 22612 22423
rect 22560 22380 22612 22389
rect 23756 22380 23808 22432
rect 25964 22380 26016 22432
rect 33324 22380 33376 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 17132 22176 17184 22228
rect 12440 22108 12492 22160
rect 19524 22176 19576 22228
rect 19984 22176 20036 22228
rect 21272 22176 21324 22228
rect 24400 22176 24452 22228
rect 25596 22176 25648 22228
rect 25964 22176 26016 22228
rect 27804 22219 27856 22228
rect 27804 22185 27813 22219
rect 27813 22185 27847 22219
rect 27847 22185 27856 22219
rect 27804 22176 27856 22185
rect 28448 22176 28500 22228
rect 29644 22219 29696 22228
rect 29644 22185 29653 22219
rect 29653 22185 29687 22219
rect 29687 22185 29696 22219
rect 29644 22176 29696 22185
rect 30380 22176 30432 22228
rect 33324 22176 33376 22228
rect 13084 21972 13136 22024
rect 14464 22040 14516 22092
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 15292 21972 15344 22024
rect 19340 22108 19392 22160
rect 20168 22108 20220 22160
rect 16764 22040 16816 22092
rect 15568 21972 15620 22024
rect 16212 22015 16264 22024
rect 14280 21904 14332 21956
rect 13452 21836 13504 21888
rect 15108 21947 15160 21956
rect 15108 21913 15117 21947
rect 15117 21913 15151 21947
rect 15151 21913 15160 21947
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 18144 22040 18196 22092
rect 20904 22083 20956 22092
rect 20904 22049 20913 22083
rect 20913 22049 20947 22083
rect 20947 22049 20956 22083
rect 20904 22040 20956 22049
rect 24584 22040 24636 22092
rect 26976 22108 27028 22160
rect 29552 22108 29604 22160
rect 25504 22083 25556 22092
rect 17316 21947 17368 21956
rect 15108 21904 15160 21913
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 17316 21913 17325 21947
rect 17325 21913 17359 21947
rect 17359 21913 17368 21947
rect 17316 21904 17368 21913
rect 15384 21836 15436 21845
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 16488 21836 16540 21888
rect 18236 21972 18288 22024
rect 19340 21972 19392 22024
rect 20536 21972 20588 22024
rect 20628 22015 20680 22024
rect 20628 21981 20637 22015
rect 20637 21981 20671 22015
rect 20671 21981 20680 22015
rect 20628 21972 20680 21981
rect 23112 21972 23164 22024
rect 24860 21972 24912 22024
rect 19984 21836 20036 21888
rect 23020 21904 23072 21956
rect 24216 21904 24268 21956
rect 24492 21947 24544 21956
rect 24492 21913 24501 21947
rect 24501 21913 24535 21947
rect 24535 21913 24544 21947
rect 24492 21904 24544 21913
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 25504 22049 25513 22083
rect 25513 22049 25547 22083
rect 25547 22049 25556 22083
rect 25504 22040 25556 22049
rect 28172 22040 28224 22092
rect 25872 21972 25924 22024
rect 26240 21972 26292 22024
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 27896 21972 27948 22024
rect 26332 21879 26384 21888
rect 26332 21845 26341 21879
rect 26341 21845 26375 21879
rect 26375 21845 26384 21879
rect 26332 21836 26384 21845
rect 26516 21879 26568 21888
rect 26516 21845 26525 21879
rect 26525 21845 26559 21879
rect 26559 21845 26568 21879
rect 26516 21836 26568 21845
rect 27528 21879 27580 21888
rect 27528 21845 27537 21879
rect 27537 21845 27571 21879
rect 27571 21845 27580 21879
rect 27528 21836 27580 21845
rect 28356 21972 28408 22024
rect 29920 22040 29972 22092
rect 30196 22040 30248 22092
rect 29644 21972 29696 22024
rect 30288 22015 30340 22024
rect 30288 21981 30297 22015
rect 30297 21981 30331 22015
rect 30331 21981 30340 22015
rect 30288 21972 30340 21981
rect 32496 22108 32548 22160
rect 32680 22083 32732 22092
rect 32680 22049 32689 22083
rect 32689 22049 32723 22083
rect 32723 22049 32732 22083
rect 32680 22040 32732 22049
rect 33324 22040 33376 22092
rect 34796 22040 34848 22092
rect 31300 21972 31352 22024
rect 32128 21972 32180 22024
rect 32496 21972 32548 22024
rect 33048 21972 33100 22024
rect 34704 21972 34756 22024
rect 29828 21947 29880 21956
rect 29828 21913 29837 21947
rect 29837 21913 29871 21947
rect 29871 21913 29880 21947
rect 29828 21904 29880 21913
rect 33600 21947 33652 21956
rect 33140 21879 33192 21888
rect 33140 21845 33149 21879
rect 33149 21845 33183 21879
rect 33183 21845 33192 21879
rect 33140 21836 33192 21845
rect 33600 21913 33609 21947
rect 33609 21913 33643 21947
rect 33643 21913 33652 21947
rect 33600 21904 33652 21913
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 15292 21632 15344 21684
rect 16488 21632 16540 21684
rect 17776 21632 17828 21684
rect 20168 21632 20220 21684
rect 20628 21632 20680 21684
rect 24308 21632 24360 21684
rect 25412 21632 25464 21684
rect 26056 21632 26108 21684
rect 26976 21632 27028 21684
rect 31208 21675 31260 21684
rect 15108 21564 15160 21616
rect 16304 21564 16356 21616
rect 21824 21607 21876 21616
rect 21824 21573 21833 21607
rect 21833 21573 21867 21607
rect 21867 21573 21876 21607
rect 21824 21564 21876 21573
rect 22008 21607 22060 21616
rect 22008 21573 22033 21607
rect 22033 21573 22060 21607
rect 22008 21564 22060 21573
rect 23020 21564 23072 21616
rect 25596 21607 25648 21616
rect 12808 21539 12860 21548
rect 12808 21505 12817 21539
rect 12817 21505 12851 21539
rect 12851 21505 12860 21539
rect 12808 21496 12860 21505
rect 13084 21539 13136 21548
rect 13084 21505 13118 21539
rect 13118 21505 13136 21539
rect 13084 21496 13136 21505
rect 14832 21496 14884 21548
rect 15752 21496 15804 21548
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 18144 21496 18196 21548
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 20720 21539 20772 21548
rect 20720 21505 20729 21539
rect 20729 21505 20763 21539
rect 20763 21505 20772 21539
rect 20720 21496 20772 21505
rect 13820 21428 13872 21480
rect 14280 21292 14332 21344
rect 16396 21360 16448 21412
rect 15476 21292 15528 21344
rect 17316 21292 17368 21344
rect 19248 21292 19300 21344
rect 20996 21292 21048 21344
rect 22560 21496 22612 21548
rect 25596 21573 25605 21607
rect 25605 21573 25639 21607
rect 25639 21573 25648 21607
rect 25596 21564 25648 21573
rect 25964 21564 26016 21616
rect 27988 21564 28040 21616
rect 23480 21496 23532 21548
rect 24860 21496 24912 21548
rect 25688 21496 25740 21548
rect 26516 21496 26568 21548
rect 27528 21496 27580 21548
rect 31208 21641 31217 21675
rect 31217 21641 31251 21675
rect 31251 21641 31260 21675
rect 31208 21632 31260 21641
rect 32680 21632 32732 21684
rect 33600 21632 33652 21684
rect 33140 21564 33192 21616
rect 33876 21564 33928 21616
rect 28448 21539 28500 21548
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 25964 21428 26016 21480
rect 27712 21428 27764 21480
rect 28448 21505 28457 21539
rect 28457 21505 28491 21539
rect 28491 21505 28500 21539
rect 28448 21496 28500 21505
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 29552 21539 29604 21548
rect 29552 21505 29561 21539
rect 29561 21505 29595 21539
rect 29595 21505 29604 21539
rect 29552 21496 29604 21505
rect 30012 21496 30064 21548
rect 30196 21539 30248 21548
rect 30196 21505 30205 21539
rect 30205 21505 30239 21539
rect 30239 21505 30248 21539
rect 30196 21496 30248 21505
rect 31300 21496 31352 21548
rect 32312 21539 32364 21548
rect 29644 21428 29696 21480
rect 30104 21428 30156 21480
rect 30564 21428 30616 21480
rect 23664 21360 23716 21412
rect 24768 21360 24820 21412
rect 23756 21335 23808 21344
rect 23756 21301 23765 21335
rect 23765 21301 23799 21335
rect 23799 21301 23808 21335
rect 23756 21292 23808 21301
rect 25320 21292 25372 21344
rect 26148 21292 26200 21344
rect 27804 21335 27856 21344
rect 27804 21301 27813 21335
rect 27813 21301 27847 21335
rect 27847 21301 27856 21335
rect 27804 21292 27856 21301
rect 28724 21292 28776 21344
rect 29000 21292 29052 21344
rect 29920 21292 29972 21344
rect 30288 21335 30340 21344
rect 30288 21301 30297 21335
rect 30297 21301 30331 21335
rect 30331 21301 30340 21335
rect 30288 21292 30340 21301
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32404 21496 32456 21548
rect 32312 21360 32364 21412
rect 32864 21496 32916 21548
rect 34796 21496 34848 21548
rect 33508 21471 33560 21480
rect 33508 21437 33517 21471
rect 33517 21437 33551 21471
rect 33551 21437 33560 21471
rect 33508 21428 33560 21437
rect 35624 21471 35676 21480
rect 35624 21437 35633 21471
rect 35633 21437 35667 21471
rect 35667 21437 35676 21471
rect 35624 21428 35676 21437
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13084 21088 13136 21140
rect 14832 21088 14884 21140
rect 15476 21088 15528 21140
rect 16396 21088 16448 21140
rect 19064 21088 19116 21140
rect 16580 21020 16632 21072
rect 16948 21020 17000 21072
rect 19984 21088 20036 21140
rect 21824 21088 21876 21140
rect 23756 21088 23808 21140
rect 25136 21088 25188 21140
rect 25780 21088 25832 21140
rect 22652 21063 22704 21072
rect 15108 20952 15160 21004
rect 13452 20927 13504 20936
rect 13452 20893 13461 20927
rect 13461 20893 13495 20927
rect 13495 20893 13504 20927
rect 13452 20884 13504 20893
rect 15200 20884 15252 20936
rect 15568 20884 15620 20936
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 16764 20927 16816 20936
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 16764 20884 16816 20893
rect 16028 20816 16080 20868
rect 17040 20884 17092 20936
rect 19340 20952 19392 21004
rect 22652 21029 22661 21063
rect 22661 21029 22695 21063
rect 22695 21029 22704 21063
rect 22652 21020 22704 21029
rect 22744 21020 22796 21072
rect 23204 21020 23256 21072
rect 23296 21020 23348 21072
rect 26424 21088 26476 21140
rect 27252 21088 27304 21140
rect 28264 21088 28316 21140
rect 28908 21088 28960 21140
rect 29184 21088 29236 21140
rect 29276 21088 29328 21140
rect 29920 21088 29972 21140
rect 32312 21131 32364 21140
rect 32312 21097 32321 21131
rect 32321 21097 32355 21131
rect 32355 21097 32364 21131
rect 32312 21088 32364 21097
rect 32496 21088 32548 21140
rect 27712 21020 27764 21072
rect 28816 21020 28868 21072
rect 30196 21020 30248 21072
rect 18420 20927 18472 20936
rect 18420 20893 18429 20927
rect 18429 20893 18463 20927
rect 18463 20893 18472 20927
rect 18420 20884 18472 20893
rect 19064 20884 19116 20936
rect 19156 20884 19208 20936
rect 20076 20884 20128 20936
rect 24860 20952 24912 21004
rect 26976 20952 27028 21004
rect 27896 20952 27948 21004
rect 17684 20816 17736 20868
rect 21456 20816 21508 20868
rect 18052 20791 18104 20800
rect 18052 20757 18061 20791
rect 18061 20757 18095 20791
rect 18095 20757 18104 20791
rect 18052 20748 18104 20757
rect 20536 20791 20588 20800
rect 20536 20757 20545 20791
rect 20545 20757 20579 20791
rect 20579 20757 20588 20791
rect 20536 20748 20588 20757
rect 22192 20748 22244 20800
rect 22836 20748 22888 20800
rect 23480 20884 23532 20936
rect 25320 20884 25372 20936
rect 26792 20884 26844 20936
rect 27436 20884 27488 20936
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 29092 20952 29144 21004
rect 27528 20884 27580 20893
rect 24216 20816 24268 20868
rect 25504 20816 25556 20868
rect 26240 20816 26292 20868
rect 23572 20748 23624 20800
rect 26424 20748 26476 20800
rect 28448 20816 28500 20868
rect 28632 20893 28643 20914
rect 28643 20893 28677 20914
rect 28677 20893 28684 20914
rect 28632 20862 28684 20893
rect 29000 20927 29052 20936
rect 29000 20893 29009 20927
rect 29009 20893 29043 20927
rect 29043 20893 29052 20927
rect 29000 20884 29052 20893
rect 28724 20859 28776 20868
rect 28724 20825 28733 20859
rect 28733 20825 28767 20859
rect 28767 20825 28776 20859
rect 28724 20816 28776 20825
rect 29092 20816 29144 20868
rect 29184 20816 29236 20868
rect 30564 20884 30616 20936
rect 32772 21020 32824 21072
rect 32864 21020 32916 21072
rect 32404 20995 32456 21004
rect 32404 20961 32413 20995
rect 32413 20961 32447 20995
rect 32447 20961 32456 20995
rect 32404 20952 32456 20961
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 33324 20995 33376 21004
rect 33324 20961 33333 20995
rect 33333 20961 33367 20995
rect 33367 20961 33376 20995
rect 33324 20952 33376 20961
rect 33876 20884 33928 20936
rect 29552 20748 29604 20800
rect 29828 20748 29880 20800
rect 30840 20748 30892 20800
rect 32772 20748 32824 20800
rect 33416 20791 33468 20800
rect 33416 20757 33425 20791
rect 33425 20757 33459 20791
rect 33459 20757 33468 20791
rect 33416 20748 33468 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 12808 20544 12860 20596
rect 15108 20544 15160 20596
rect 18512 20544 18564 20596
rect 21640 20544 21692 20596
rect 13452 20476 13504 20528
rect 18052 20476 18104 20528
rect 20996 20476 21048 20528
rect 22652 20544 22704 20596
rect 23204 20544 23256 20596
rect 26240 20587 26292 20596
rect 26240 20553 26249 20587
rect 26249 20553 26283 20587
rect 26283 20553 26292 20587
rect 26240 20544 26292 20553
rect 26424 20544 26476 20596
rect 28540 20544 28592 20596
rect 28632 20544 28684 20596
rect 28908 20587 28960 20596
rect 28908 20553 28917 20587
rect 28917 20553 28951 20587
rect 28951 20553 28960 20587
rect 28908 20544 28960 20553
rect 29828 20544 29880 20596
rect 32588 20544 32640 20596
rect 32772 20544 32824 20596
rect 32956 20544 33008 20596
rect 34796 20544 34848 20596
rect 12624 20408 12676 20460
rect 13728 20408 13780 20460
rect 13912 20451 13964 20460
rect 13912 20417 13946 20451
rect 13946 20417 13964 20451
rect 13912 20408 13964 20417
rect 16396 20408 16448 20460
rect 19248 20408 19300 20460
rect 21088 20408 21140 20460
rect 21640 20408 21692 20460
rect 21732 20408 21784 20460
rect 23112 20451 23164 20460
rect 23112 20417 23121 20451
rect 23121 20417 23155 20451
rect 23155 20417 23164 20451
rect 23112 20408 23164 20417
rect 23388 20451 23440 20460
rect 23388 20417 23422 20451
rect 23422 20417 23440 20451
rect 23388 20408 23440 20417
rect 24860 20408 24912 20460
rect 27252 20476 27304 20528
rect 33416 20476 33468 20528
rect 15476 20340 15528 20392
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 20444 20340 20496 20392
rect 21180 20383 21232 20392
rect 21180 20349 21189 20383
rect 21189 20349 21223 20383
rect 21223 20349 21232 20383
rect 21180 20340 21232 20349
rect 24676 20340 24728 20392
rect 25504 20340 25556 20392
rect 27804 20408 27856 20460
rect 29736 20408 29788 20460
rect 30288 20451 30340 20460
rect 30288 20417 30297 20451
rect 30297 20417 30331 20451
rect 30331 20417 30340 20451
rect 30288 20408 30340 20417
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 33324 20408 33376 20460
rect 33508 20451 33560 20460
rect 33508 20417 33517 20451
rect 33517 20417 33551 20451
rect 33551 20417 33560 20451
rect 33508 20408 33560 20417
rect 19064 20272 19116 20324
rect 25596 20272 25648 20324
rect 27344 20272 27396 20324
rect 15568 20204 15620 20256
rect 21180 20204 21232 20256
rect 23112 20204 23164 20256
rect 24308 20204 24360 20256
rect 28540 20340 28592 20392
rect 28724 20383 28776 20392
rect 28724 20349 28733 20383
rect 28733 20349 28767 20383
rect 28767 20349 28776 20383
rect 28724 20340 28776 20349
rect 28080 20272 28132 20324
rect 30472 20383 30524 20392
rect 30472 20349 30481 20383
rect 30481 20349 30515 20383
rect 30515 20349 30524 20383
rect 30472 20340 30524 20349
rect 29920 20315 29972 20324
rect 28172 20204 28224 20256
rect 28724 20204 28776 20256
rect 29920 20281 29929 20315
rect 29929 20281 29963 20315
rect 29963 20281 29972 20315
rect 29920 20272 29972 20281
rect 30288 20272 30340 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 13912 20000 13964 20052
rect 20536 20000 20588 20052
rect 17316 19932 17368 19984
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 15384 19864 15436 19916
rect 17040 19864 17092 19916
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 15568 19796 15620 19848
rect 16212 19796 16264 19848
rect 16948 19796 17000 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 20720 19932 20772 19984
rect 21456 20000 21508 20052
rect 23388 20043 23440 20052
rect 23388 20009 23397 20043
rect 23397 20009 23431 20043
rect 23431 20009 23440 20043
rect 23388 20000 23440 20009
rect 22100 19932 22152 19984
rect 22192 19932 22244 19984
rect 24584 20000 24636 20052
rect 27528 20000 27580 20052
rect 30564 20043 30616 20052
rect 24492 19932 24544 19984
rect 25136 19932 25188 19984
rect 28080 19932 28132 19984
rect 30564 20009 30573 20043
rect 30573 20009 30607 20043
rect 30607 20009 30616 20043
rect 30564 20000 30616 20009
rect 32864 20000 32916 20052
rect 35348 19975 35400 19984
rect 17776 19796 17828 19805
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 20260 19839 20312 19848
rect 16396 19728 16448 19780
rect 16948 19660 17000 19712
rect 18788 19728 18840 19780
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20628 19796 20680 19848
rect 20720 19728 20772 19780
rect 18328 19660 18380 19712
rect 21180 19660 21232 19712
rect 21272 19660 21324 19712
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 22100 19839 22152 19848
rect 21456 19796 21508 19805
rect 22100 19805 22109 19839
rect 22109 19805 22143 19839
rect 22143 19805 22152 19839
rect 22100 19796 22152 19805
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 23480 19796 23532 19848
rect 24860 19796 24912 19848
rect 24676 19728 24728 19780
rect 25780 19796 25832 19848
rect 26516 19796 26568 19848
rect 29552 19796 29604 19848
rect 30472 19796 30524 19848
rect 27252 19771 27304 19780
rect 21456 19660 21508 19712
rect 21824 19660 21876 19712
rect 23480 19660 23532 19712
rect 24308 19660 24360 19712
rect 27252 19737 27261 19771
rect 27261 19737 27295 19771
rect 27295 19737 27304 19771
rect 27252 19728 27304 19737
rect 28264 19771 28316 19780
rect 28264 19737 28273 19771
rect 28273 19737 28307 19771
rect 28307 19737 28316 19771
rect 28264 19728 28316 19737
rect 28816 19728 28868 19780
rect 31392 19864 31444 19916
rect 33140 19864 33192 19916
rect 30656 19796 30708 19848
rect 30932 19839 30984 19848
rect 30932 19805 30941 19839
rect 30941 19805 30975 19839
rect 30975 19805 30984 19839
rect 30932 19796 30984 19805
rect 31024 19796 31076 19848
rect 32588 19796 32640 19848
rect 33048 19796 33100 19848
rect 33416 19796 33468 19848
rect 35348 19941 35357 19975
rect 35357 19941 35391 19975
rect 35391 19941 35400 19975
rect 35348 19932 35400 19941
rect 25320 19660 25372 19712
rect 28448 19660 28500 19712
rect 33784 19728 33836 19780
rect 32956 19660 33008 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 20260 19456 20312 19508
rect 13452 19431 13504 19440
rect 13452 19397 13461 19431
rect 13461 19397 13495 19431
rect 13495 19397 13504 19431
rect 13452 19388 13504 19397
rect 17132 19388 17184 19440
rect 19248 19388 19300 19440
rect 20996 19456 21048 19508
rect 22192 19456 22244 19508
rect 25044 19456 25096 19508
rect 27252 19456 27304 19508
rect 27436 19499 27488 19508
rect 27436 19465 27445 19499
rect 27445 19465 27479 19499
rect 27479 19465 27488 19499
rect 27436 19456 27488 19465
rect 28080 19499 28132 19508
rect 28080 19465 28089 19499
rect 28089 19465 28123 19499
rect 28123 19465 28132 19499
rect 28080 19456 28132 19465
rect 32312 19456 32364 19508
rect 32956 19499 33008 19508
rect 32956 19465 32965 19499
rect 32965 19465 32999 19499
rect 32999 19465 33008 19499
rect 32956 19456 33008 19465
rect 33784 19499 33836 19508
rect 33784 19465 33793 19499
rect 33793 19465 33827 19499
rect 33827 19465 33836 19499
rect 33784 19456 33836 19465
rect 11888 19320 11940 19372
rect 15384 19320 15436 19372
rect 16856 19363 16908 19372
rect 15108 19184 15160 19236
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 18328 19363 18380 19372
rect 18328 19329 18337 19363
rect 18337 19329 18371 19363
rect 18371 19329 18380 19363
rect 18328 19320 18380 19329
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 18788 19320 18840 19372
rect 21824 19388 21876 19440
rect 24492 19388 24544 19440
rect 16764 19252 16816 19304
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 19156 19252 19208 19304
rect 17224 19184 17276 19236
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20536 19363 20588 19372
rect 20076 19320 20128 19329
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20812 19363 20864 19372
rect 20260 19252 20312 19304
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 12624 19116 12676 19168
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 16580 19116 16632 19168
rect 20076 19116 20128 19168
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 20996 19320 21048 19372
rect 21548 19320 21600 19372
rect 22836 19363 22888 19372
rect 22836 19329 22870 19363
rect 22870 19329 22888 19363
rect 22836 19320 22888 19329
rect 23572 19320 23624 19372
rect 24768 19320 24820 19372
rect 25412 19363 25464 19372
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 25872 19252 25924 19304
rect 27528 19363 27580 19372
rect 27528 19329 27537 19363
rect 27537 19329 27571 19363
rect 27571 19329 27580 19363
rect 27528 19320 27580 19329
rect 28816 19388 28868 19440
rect 30380 19388 30432 19440
rect 30932 19388 30984 19440
rect 32864 19431 32916 19440
rect 32864 19397 32873 19431
rect 32873 19397 32907 19431
rect 32907 19397 32916 19431
rect 32864 19388 32916 19397
rect 34796 19388 34848 19440
rect 29368 19363 29420 19372
rect 23756 19116 23808 19168
rect 24032 19116 24084 19168
rect 27620 19295 27672 19304
rect 27620 19261 27629 19295
rect 27629 19261 27663 19295
rect 27663 19261 27672 19295
rect 27620 19252 27672 19261
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 29552 19363 29604 19372
rect 29552 19329 29561 19363
rect 29561 19329 29595 19363
rect 29595 19329 29604 19363
rect 29552 19320 29604 19329
rect 30840 19363 30892 19372
rect 30840 19329 30849 19363
rect 30849 19329 30883 19363
rect 30883 19329 30892 19363
rect 30840 19320 30892 19329
rect 32404 19320 32456 19372
rect 29644 19295 29696 19304
rect 29644 19261 29653 19295
rect 29653 19261 29687 19295
rect 29687 19261 29696 19295
rect 29644 19252 29696 19261
rect 33140 19295 33192 19304
rect 33140 19261 33149 19295
rect 33149 19261 33183 19295
rect 33183 19261 33192 19295
rect 33140 19252 33192 19261
rect 28632 19184 28684 19236
rect 30380 19227 30432 19236
rect 30380 19193 30389 19227
rect 30389 19193 30423 19227
rect 30423 19193 30432 19227
rect 30380 19184 30432 19193
rect 29184 19159 29236 19168
rect 29184 19125 29193 19159
rect 29193 19125 29227 19159
rect 29227 19125 29236 19159
rect 29184 19116 29236 19125
rect 29736 19116 29788 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 13452 18955 13504 18964
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 16396 18955 16448 18964
rect 16396 18921 16405 18955
rect 16405 18921 16439 18955
rect 16439 18921 16448 18955
rect 16396 18912 16448 18921
rect 19892 18912 19944 18964
rect 15476 18844 15528 18896
rect 20904 18912 20956 18964
rect 22100 18912 22152 18964
rect 23296 18955 23348 18964
rect 23296 18921 23305 18955
rect 23305 18921 23339 18955
rect 23339 18921 23348 18955
rect 23296 18912 23348 18921
rect 20720 18844 20772 18896
rect 16948 18776 17000 18828
rect 17316 18776 17368 18828
rect 17868 18819 17920 18828
rect 17868 18785 17877 18819
rect 17877 18785 17911 18819
rect 17911 18785 17920 18819
rect 17868 18776 17920 18785
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 12808 18708 12860 18760
rect 13728 18708 13780 18760
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 11060 18640 11112 18692
rect 13360 18683 13412 18692
rect 13360 18649 13369 18683
rect 13369 18649 13403 18683
rect 13403 18649 13412 18683
rect 13360 18640 13412 18649
rect 13820 18640 13872 18692
rect 15936 18640 15988 18692
rect 17224 18708 17276 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 18604 18708 18656 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 18512 18640 18564 18692
rect 19340 18640 19392 18692
rect 11796 18572 11848 18624
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 16856 18572 16908 18624
rect 17684 18572 17736 18624
rect 19432 18572 19484 18624
rect 21088 18776 21140 18828
rect 21548 18776 21600 18828
rect 26240 18912 26292 18964
rect 27620 18912 27672 18964
rect 29644 18912 29696 18964
rect 30288 18912 30340 18964
rect 32220 18912 32272 18964
rect 33324 18912 33376 18964
rect 23572 18887 23624 18896
rect 23572 18853 23581 18887
rect 23581 18853 23615 18887
rect 23615 18853 23624 18887
rect 23572 18844 23624 18853
rect 23664 18887 23716 18896
rect 23664 18853 23673 18887
rect 23673 18853 23707 18887
rect 23707 18853 23716 18887
rect 23664 18844 23716 18853
rect 25228 18844 25280 18896
rect 19984 18708 20036 18760
rect 19800 18683 19852 18692
rect 19800 18649 19809 18683
rect 19809 18649 19843 18683
rect 19843 18649 19852 18683
rect 19800 18640 19852 18649
rect 20628 18751 20680 18760
rect 20628 18717 20638 18751
rect 20638 18717 20672 18751
rect 20672 18717 20680 18751
rect 20628 18708 20680 18717
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 20996 18751 21048 18760
rect 20996 18717 21010 18751
rect 21010 18717 21044 18751
rect 21044 18717 21048 18751
rect 21640 18751 21692 18760
rect 20996 18708 21048 18717
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 22468 18708 22520 18760
rect 24032 18776 24084 18828
rect 25320 18819 25372 18828
rect 25320 18785 25329 18819
rect 25329 18785 25363 18819
rect 25363 18785 25372 18819
rect 25320 18776 25372 18785
rect 27160 18776 27212 18828
rect 29460 18844 29512 18896
rect 32772 18844 32824 18896
rect 27988 18776 28040 18828
rect 29092 18776 29144 18828
rect 23756 18751 23808 18760
rect 23756 18717 23765 18751
rect 23765 18717 23799 18751
rect 23799 18717 23808 18751
rect 23756 18708 23808 18717
rect 20812 18572 20864 18624
rect 22928 18640 22980 18692
rect 23204 18640 23256 18692
rect 24584 18683 24636 18692
rect 24584 18649 24593 18683
rect 24593 18649 24627 18683
rect 24627 18649 24636 18683
rect 24584 18640 24636 18649
rect 25872 18640 25924 18692
rect 27712 18751 27764 18760
rect 27712 18717 27721 18751
rect 27721 18717 27755 18751
rect 27755 18717 27764 18751
rect 27712 18708 27764 18717
rect 28080 18708 28132 18760
rect 28356 18708 28408 18760
rect 28724 18751 28776 18760
rect 28724 18717 28733 18751
rect 28733 18717 28767 18751
rect 28767 18717 28776 18751
rect 28724 18708 28776 18717
rect 29276 18708 29328 18760
rect 30196 18751 30248 18760
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 30196 18708 30248 18717
rect 30472 18751 30524 18760
rect 28172 18640 28224 18692
rect 30104 18640 30156 18692
rect 30472 18717 30481 18751
rect 30481 18717 30515 18751
rect 30515 18717 30524 18751
rect 30472 18708 30524 18717
rect 30564 18751 30616 18760
rect 30564 18717 30573 18751
rect 30573 18717 30607 18751
rect 30607 18717 30616 18751
rect 30564 18708 30616 18717
rect 32036 18708 32088 18760
rect 33232 18776 33284 18828
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 32956 18683 33008 18692
rect 32956 18649 32965 18683
rect 32965 18649 32999 18683
rect 32999 18649 33008 18683
rect 32956 18640 33008 18649
rect 22192 18572 22244 18624
rect 23112 18572 23164 18624
rect 24860 18572 24912 18624
rect 25320 18572 25372 18624
rect 26608 18572 26660 18624
rect 27160 18572 27212 18624
rect 29000 18615 29052 18624
rect 29000 18581 29009 18615
rect 29009 18581 29043 18615
rect 29043 18581 29052 18615
rect 29000 18572 29052 18581
rect 32588 18572 32640 18624
rect 33324 18615 33376 18624
rect 33324 18581 33333 18615
rect 33333 18581 33367 18615
rect 33367 18581 33376 18615
rect 33324 18572 33376 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 15016 18368 15068 18420
rect 19984 18368 20036 18420
rect 21272 18411 21324 18420
rect 10692 18232 10744 18284
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 14556 18232 14608 18284
rect 18144 18300 18196 18352
rect 19524 18300 19576 18352
rect 15936 18232 15988 18284
rect 16212 18232 16264 18284
rect 19248 18232 19300 18284
rect 11520 18207 11572 18216
rect 11520 18173 11529 18207
rect 11529 18173 11563 18207
rect 11563 18173 11572 18207
rect 11520 18164 11572 18173
rect 12532 18028 12584 18080
rect 14464 18028 14516 18080
rect 15568 18028 15620 18080
rect 15752 18028 15804 18080
rect 17040 18164 17092 18216
rect 19064 18164 19116 18216
rect 17960 18096 18012 18148
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 22284 18368 22336 18420
rect 22468 18368 22520 18420
rect 20904 18232 20956 18241
rect 22008 18232 22060 18284
rect 23020 18368 23072 18420
rect 17040 18028 17092 18080
rect 19524 18028 19576 18080
rect 19616 18028 19668 18080
rect 20720 18096 20772 18148
rect 21272 18164 21324 18216
rect 22928 18232 22980 18284
rect 25596 18368 25648 18420
rect 28080 18368 28132 18420
rect 29368 18368 29420 18420
rect 30564 18368 30616 18420
rect 30656 18368 30708 18420
rect 32496 18368 32548 18420
rect 33600 18368 33652 18420
rect 25228 18300 25280 18352
rect 28264 18300 28316 18352
rect 31024 18343 31076 18352
rect 31024 18309 31033 18343
rect 31033 18309 31067 18343
rect 31067 18309 31076 18343
rect 31024 18300 31076 18309
rect 32404 18300 32456 18352
rect 33692 18300 33744 18352
rect 33876 18300 33928 18352
rect 22652 18164 22704 18216
rect 22836 18164 22888 18216
rect 23020 18164 23072 18216
rect 23204 18164 23256 18216
rect 24492 18275 24544 18284
rect 24492 18241 24501 18275
rect 24501 18241 24535 18275
rect 24535 18241 24544 18275
rect 24492 18232 24544 18241
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 25320 18275 25372 18284
rect 24676 18232 24728 18241
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 25872 18232 25924 18284
rect 20904 18096 20956 18148
rect 24584 18096 24636 18148
rect 24860 18096 24912 18148
rect 25504 18096 25556 18148
rect 27068 18232 27120 18284
rect 27804 18232 27856 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 28724 18232 28776 18284
rect 29092 18232 29144 18284
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 28264 18207 28316 18216
rect 28264 18173 28273 18207
rect 28273 18173 28307 18207
rect 28307 18173 28316 18207
rect 28264 18164 28316 18173
rect 29276 18164 29328 18216
rect 30288 18232 30340 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 32588 18232 32640 18284
rect 30104 18164 30156 18216
rect 32864 18164 32916 18216
rect 33232 18232 33284 18284
rect 33600 18232 33652 18284
rect 34152 18281 34204 18284
rect 34152 18247 34166 18281
rect 34166 18247 34200 18281
rect 34200 18247 34204 18281
rect 34152 18232 34204 18247
rect 27620 18096 27672 18148
rect 28908 18096 28960 18148
rect 30932 18096 30984 18148
rect 31392 18096 31444 18148
rect 22376 18028 22428 18080
rect 23020 18071 23072 18080
rect 23020 18037 23029 18071
rect 23029 18037 23063 18071
rect 23063 18037 23072 18071
rect 23020 18028 23072 18037
rect 23388 18071 23440 18080
rect 23388 18037 23397 18071
rect 23397 18037 23431 18071
rect 23431 18037 23440 18071
rect 23388 18028 23440 18037
rect 24952 18028 25004 18080
rect 27528 18028 27580 18080
rect 29368 18028 29420 18080
rect 31760 18028 31812 18080
rect 32956 18028 33008 18080
rect 33140 18028 33192 18080
rect 34152 18028 34204 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 11796 17824 11848 17876
rect 14556 17867 14608 17876
rect 14556 17833 14565 17867
rect 14565 17833 14599 17867
rect 14599 17833 14608 17867
rect 14556 17824 14608 17833
rect 16856 17824 16908 17876
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 18144 17824 18196 17876
rect 19248 17867 19300 17876
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 21180 17867 21232 17876
rect 21180 17833 21189 17867
rect 21189 17833 21223 17867
rect 21223 17833 21232 17867
rect 21180 17824 21232 17833
rect 11428 17731 11480 17740
rect 11428 17697 11437 17731
rect 11437 17697 11471 17731
rect 11471 17697 11480 17731
rect 11428 17688 11480 17697
rect 18512 17756 18564 17808
rect 20812 17756 20864 17808
rect 28080 17824 28132 17876
rect 29184 17824 29236 17876
rect 29644 17824 29696 17876
rect 23112 17756 23164 17808
rect 27804 17756 27856 17808
rect 33324 17824 33376 17876
rect 15016 17731 15068 17740
rect 15016 17697 15025 17731
rect 15025 17697 15059 17731
rect 15059 17697 15068 17731
rect 15016 17688 15068 17697
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 19524 17688 19576 17740
rect 12072 17620 12124 17672
rect 14556 17620 14608 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15108 17620 15160 17672
rect 10600 17595 10652 17604
rect 10600 17561 10609 17595
rect 10609 17561 10643 17595
rect 10643 17561 10652 17595
rect 10600 17552 10652 17561
rect 11612 17552 11664 17604
rect 13728 17552 13780 17604
rect 15384 17552 15436 17604
rect 15752 17620 15804 17672
rect 17224 17620 17276 17672
rect 17684 17663 17736 17672
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 16212 17552 16264 17604
rect 10968 17527 11020 17536
rect 10968 17493 10977 17527
rect 10977 17493 11011 17527
rect 11011 17493 11020 17527
rect 10968 17484 11020 17493
rect 11704 17484 11756 17536
rect 14556 17484 14608 17536
rect 17224 17484 17276 17536
rect 17500 17484 17552 17536
rect 18880 17620 18932 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 20076 17620 20128 17672
rect 20536 17663 20588 17672
rect 20536 17629 20545 17663
rect 20545 17629 20579 17663
rect 20579 17629 20588 17663
rect 20536 17620 20588 17629
rect 20720 17620 20772 17672
rect 22468 17688 22520 17740
rect 20996 17663 21048 17672
rect 20996 17629 21010 17663
rect 21010 17629 21044 17663
rect 21044 17629 21048 17663
rect 22928 17663 22980 17672
rect 20996 17620 21048 17629
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 23204 17688 23256 17740
rect 26792 17731 26844 17740
rect 26792 17697 26801 17731
rect 26801 17697 26835 17731
rect 26835 17697 26844 17731
rect 26792 17688 26844 17697
rect 30472 17756 30524 17808
rect 32036 17756 32088 17808
rect 31760 17731 31812 17740
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 23572 17620 23624 17672
rect 24860 17663 24912 17672
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 24952 17620 25004 17672
rect 29368 17620 29420 17672
rect 31760 17697 31769 17731
rect 31769 17697 31803 17731
rect 31803 17697 31812 17731
rect 31760 17688 31812 17697
rect 21180 17552 21232 17604
rect 21640 17552 21692 17604
rect 21088 17484 21140 17536
rect 24584 17552 24636 17604
rect 25596 17552 25648 17604
rect 26056 17552 26108 17604
rect 29092 17552 29144 17604
rect 30932 17620 30984 17672
rect 31392 17663 31444 17672
rect 31392 17629 31401 17663
rect 31401 17629 31435 17663
rect 31435 17629 31444 17663
rect 31392 17620 31444 17629
rect 31024 17552 31076 17604
rect 32220 17731 32272 17740
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 33416 17688 33468 17740
rect 32404 17663 32456 17672
rect 32404 17629 32413 17663
rect 32413 17629 32447 17663
rect 32447 17629 32456 17663
rect 32404 17620 32456 17629
rect 32496 17663 32548 17672
rect 32496 17629 32505 17663
rect 32505 17629 32539 17663
rect 32539 17629 32548 17663
rect 32772 17663 32824 17672
rect 32496 17620 32548 17629
rect 32772 17629 32781 17663
rect 32781 17629 32815 17663
rect 32815 17629 32824 17663
rect 32772 17620 32824 17629
rect 33600 17663 33652 17672
rect 33600 17629 33614 17663
rect 33614 17629 33648 17663
rect 33648 17629 33652 17663
rect 33600 17620 33652 17629
rect 33416 17595 33468 17604
rect 33416 17561 33425 17595
rect 33425 17561 33459 17595
rect 33459 17561 33468 17595
rect 33416 17552 33468 17561
rect 22652 17527 22704 17536
rect 22652 17493 22661 17527
rect 22661 17493 22695 17527
rect 22695 17493 22704 17527
rect 22652 17484 22704 17493
rect 24768 17484 24820 17536
rect 25872 17484 25924 17536
rect 29460 17484 29512 17536
rect 32220 17484 32272 17536
rect 32864 17484 32916 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 10600 17212 10652 17264
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 11612 17212 11664 17264
rect 12992 17280 13044 17332
rect 13820 17280 13872 17332
rect 12900 17212 12952 17264
rect 14464 17280 14516 17332
rect 14740 17280 14792 17332
rect 24584 17323 24636 17332
rect 14372 17212 14424 17264
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 14004 17144 14056 17196
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 14832 17212 14884 17264
rect 15016 17144 15068 17196
rect 11060 17008 11112 17060
rect 11244 17008 11296 17060
rect 14648 17076 14700 17128
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 19432 17212 19484 17264
rect 20628 17212 20680 17264
rect 21272 17212 21324 17264
rect 22192 17212 22244 17264
rect 22652 17212 22704 17264
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 16028 17144 16080 17196
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 19524 17187 19576 17196
rect 14924 17076 14976 17085
rect 16764 17076 16816 17128
rect 15476 17008 15528 17060
rect 16212 17008 16264 17060
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 19984 17144 20036 17196
rect 24584 17289 24593 17323
rect 24593 17289 24627 17323
rect 24627 17289 24636 17323
rect 24584 17280 24636 17289
rect 24676 17280 24728 17332
rect 23204 17212 23256 17264
rect 24492 17144 24544 17196
rect 24768 17144 24820 17196
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25412 17280 25464 17332
rect 26056 17280 26108 17332
rect 28172 17280 28224 17332
rect 29552 17280 29604 17332
rect 30472 17280 30524 17332
rect 30840 17280 30892 17332
rect 31024 17280 31076 17332
rect 32588 17323 32640 17332
rect 32588 17289 32597 17323
rect 32597 17289 32631 17323
rect 32631 17289 32640 17323
rect 32588 17280 32640 17289
rect 33600 17280 33652 17332
rect 25044 17144 25096 17153
rect 25412 17144 25464 17196
rect 19156 17076 19208 17128
rect 21732 17076 21784 17128
rect 22284 17119 22336 17128
rect 22284 17085 22293 17119
rect 22293 17085 22327 17119
rect 22327 17085 22336 17119
rect 22284 17076 22336 17085
rect 22652 17076 22704 17128
rect 25320 17076 25372 17128
rect 29000 17144 29052 17196
rect 27896 17076 27948 17128
rect 21548 17008 21600 17060
rect 24308 17008 24360 17060
rect 27436 17008 27488 17060
rect 27712 17008 27764 17060
rect 28724 17076 28776 17128
rect 31024 17144 31076 17196
rect 31668 17144 31720 17196
rect 32220 17187 32272 17196
rect 32220 17153 32229 17187
rect 32229 17153 32263 17187
rect 32263 17153 32272 17187
rect 32220 17144 32272 17153
rect 29184 17008 29236 17060
rect 29276 17008 29328 17060
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 15108 16940 15160 16992
rect 17132 16940 17184 16992
rect 19248 16940 19300 16992
rect 20536 16940 20588 16992
rect 20628 16940 20680 16992
rect 20904 16940 20956 16992
rect 21916 16940 21968 16992
rect 22928 16940 22980 16992
rect 24032 16940 24084 16992
rect 27068 16983 27120 16992
rect 27068 16949 27077 16983
rect 27077 16949 27111 16983
rect 27111 16949 27120 16983
rect 27068 16940 27120 16949
rect 28448 16940 28500 16992
rect 30840 17008 30892 17060
rect 33324 17144 33376 17196
rect 32220 16940 32272 16992
rect 33048 16940 33100 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 13728 16736 13780 16788
rect 13820 16736 13872 16788
rect 16948 16736 17000 16788
rect 19984 16779 20036 16788
rect 19984 16745 19993 16779
rect 19993 16745 20027 16779
rect 20027 16745 20036 16779
rect 19984 16736 20036 16745
rect 20536 16736 20588 16788
rect 23664 16736 23716 16788
rect 24860 16736 24912 16788
rect 11520 16643 11572 16652
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 12164 16600 12216 16652
rect 11244 16532 11296 16584
rect 12624 16532 12676 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 15752 16668 15804 16720
rect 19156 16668 19208 16720
rect 20076 16668 20128 16720
rect 23388 16668 23440 16720
rect 14188 16600 14240 16652
rect 12992 16532 13044 16541
rect 14004 16532 14056 16584
rect 14372 16532 14424 16584
rect 14740 16532 14792 16584
rect 13084 16464 13136 16516
rect 13176 16464 13228 16516
rect 10692 16396 10744 16448
rect 13452 16396 13504 16448
rect 17132 16600 17184 16652
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 15752 16532 15804 16584
rect 17592 16532 17644 16584
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 18144 16532 18196 16584
rect 18604 16600 18656 16652
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 21456 16600 21508 16652
rect 16948 16464 17000 16516
rect 17408 16464 17460 16516
rect 18788 16532 18840 16584
rect 17132 16396 17184 16448
rect 17592 16396 17644 16448
rect 19156 16464 19208 16516
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 20444 16532 20496 16584
rect 20996 16507 21048 16516
rect 20996 16473 21005 16507
rect 21005 16473 21039 16507
rect 21039 16473 21048 16507
rect 21548 16532 21600 16584
rect 22928 16532 22980 16584
rect 24308 16600 24360 16652
rect 23204 16575 23256 16584
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 23204 16532 23256 16541
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 23572 16532 23624 16584
rect 25780 16668 25832 16720
rect 25688 16600 25740 16652
rect 26792 16736 26844 16788
rect 29552 16736 29604 16788
rect 30472 16736 30524 16788
rect 33416 16736 33468 16788
rect 27436 16668 27488 16720
rect 29184 16668 29236 16720
rect 30840 16668 30892 16720
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 25596 16532 25648 16584
rect 20996 16464 21048 16473
rect 27804 16532 27856 16584
rect 29736 16600 29788 16652
rect 32220 16600 32272 16652
rect 30380 16532 30432 16584
rect 28356 16464 28408 16516
rect 30472 16464 30524 16516
rect 31668 16532 31720 16584
rect 33140 16600 33192 16652
rect 32956 16575 33008 16584
rect 21364 16396 21416 16448
rect 25596 16396 25648 16448
rect 28172 16396 28224 16448
rect 32128 16396 32180 16448
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 32956 16532 33008 16541
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 13084 16192 13136 16244
rect 13452 16124 13504 16176
rect 13544 16167 13596 16176
rect 13544 16133 13569 16167
rect 13569 16133 13596 16167
rect 15660 16192 15712 16244
rect 16764 16192 16816 16244
rect 17868 16192 17920 16244
rect 19156 16192 19208 16244
rect 21548 16192 21600 16244
rect 13544 16124 13596 16133
rect 14556 16124 14608 16176
rect 11704 16056 11756 16108
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 13636 15988 13688 16040
rect 14372 15988 14424 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 14280 15920 14332 15972
rect 15936 16056 15988 16108
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16764 16056 16816 16108
rect 17960 16124 18012 16176
rect 19708 16124 19760 16176
rect 23296 16192 23348 16244
rect 25228 16192 25280 16244
rect 30288 16235 30340 16244
rect 30288 16201 30297 16235
rect 30297 16201 30331 16235
rect 30331 16201 30340 16235
rect 30288 16192 30340 16201
rect 32404 16192 32456 16244
rect 33324 16235 33376 16244
rect 33324 16201 33333 16235
rect 33333 16201 33367 16235
rect 33367 16201 33376 16235
rect 33324 16192 33376 16201
rect 17684 16056 17736 16108
rect 18604 16099 18656 16108
rect 18236 15988 18288 16040
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 19892 16056 19944 16108
rect 20076 16099 20128 16108
rect 20076 16065 20110 16099
rect 20110 16065 20128 16099
rect 20076 16056 20128 16065
rect 21640 16056 21692 16108
rect 19616 15988 19668 16040
rect 15108 15920 15160 15972
rect 19800 15920 19852 15972
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 12256 15852 12308 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 15292 15852 15344 15904
rect 15752 15852 15804 15904
rect 18236 15852 18288 15904
rect 20996 15920 21048 15972
rect 22652 16056 22704 16108
rect 24860 16124 24912 16176
rect 24952 16124 25004 16176
rect 24400 16099 24452 16108
rect 24400 16065 24434 16099
rect 24434 16065 24452 16099
rect 24400 16056 24452 16065
rect 22008 15920 22060 15972
rect 23204 15988 23256 16040
rect 20812 15852 20864 15904
rect 21916 15852 21968 15904
rect 22192 15852 22244 15904
rect 23572 15920 23624 15972
rect 26976 16056 27028 16108
rect 27712 16056 27764 16108
rect 27988 16099 28040 16108
rect 27988 16065 27997 16099
rect 27997 16065 28031 16099
rect 28031 16065 28040 16099
rect 27988 16056 28040 16065
rect 27896 15988 27948 16040
rect 28172 16099 28224 16108
rect 28172 16065 28181 16099
rect 28181 16065 28215 16099
rect 28215 16065 28224 16099
rect 28356 16099 28408 16108
rect 28172 16056 28224 16065
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 28448 16056 28500 16108
rect 31208 16056 31260 16108
rect 32128 16099 32180 16108
rect 30656 15988 30708 16040
rect 31024 16031 31076 16040
rect 31024 15997 31033 16031
rect 31033 15997 31067 16031
rect 31067 15997 31076 16031
rect 32128 16065 32137 16099
rect 32137 16065 32171 16099
rect 32171 16065 32180 16099
rect 32128 16056 32180 16065
rect 31024 15988 31076 15997
rect 31668 15988 31720 16040
rect 28540 15920 28592 15972
rect 28724 15920 28776 15972
rect 25412 15852 25464 15904
rect 28816 15852 28868 15904
rect 28908 15895 28960 15904
rect 28908 15861 28917 15895
rect 28917 15861 28951 15895
rect 28951 15861 28960 15895
rect 30472 15920 30524 15972
rect 28908 15852 28960 15861
rect 32956 15852 33008 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 16488 15648 16540 15700
rect 24400 15691 24452 15700
rect 24400 15657 24409 15691
rect 24409 15657 24443 15691
rect 24443 15657 24452 15691
rect 24400 15648 24452 15657
rect 11796 15580 11848 15632
rect 14832 15580 14884 15632
rect 10508 15512 10560 15564
rect 14372 15512 14424 15564
rect 16396 15580 16448 15632
rect 16580 15580 16632 15632
rect 9496 15487 9548 15496
rect 9496 15453 9505 15487
rect 9505 15453 9539 15487
rect 9539 15453 9548 15487
rect 12164 15487 12216 15496
rect 9496 15444 9548 15453
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 12256 15444 12308 15496
rect 14464 15444 14516 15496
rect 15936 15512 15988 15564
rect 16764 15512 16816 15564
rect 16948 15512 17000 15564
rect 20260 15580 20312 15632
rect 11336 15419 11388 15428
rect 9680 15308 9732 15360
rect 11336 15385 11345 15419
rect 11345 15385 11379 15419
rect 11379 15385 11388 15419
rect 11336 15376 11388 15385
rect 15844 15444 15896 15496
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 16672 15444 16724 15496
rect 17960 15512 18012 15564
rect 19248 15555 19300 15564
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 19800 15512 19852 15564
rect 20996 15512 21048 15564
rect 21824 15580 21876 15632
rect 22836 15580 22888 15632
rect 24768 15580 24820 15632
rect 18144 15444 18196 15496
rect 18512 15444 18564 15496
rect 20260 15444 20312 15496
rect 21456 15444 21508 15496
rect 21824 15444 21876 15496
rect 24584 15512 24636 15564
rect 24676 15487 24728 15496
rect 24676 15453 24685 15487
rect 24685 15453 24719 15487
rect 24719 15453 24728 15487
rect 24676 15444 24728 15453
rect 27068 15648 27120 15700
rect 30472 15648 30524 15700
rect 25044 15580 25096 15632
rect 26884 15623 26936 15632
rect 26884 15589 26893 15623
rect 26893 15589 26927 15623
rect 26927 15589 26936 15623
rect 26884 15580 26936 15589
rect 28356 15512 28408 15564
rect 25320 15444 25372 15496
rect 25596 15444 25648 15496
rect 10968 15308 11020 15360
rect 15200 15308 15252 15360
rect 17132 15376 17184 15428
rect 20720 15376 20772 15428
rect 16580 15308 16632 15360
rect 16856 15308 16908 15360
rect 17500 15308 17552 15360
rect 22468 15308 22520 15360
rect 24584 15308 24636 15360
rect 27896 15376 27948 15428
rect 28264 15487 28316 15496
rect 28264 15453 28273 15487
rect 28273 15453 28307 15487
rect 28307 15453 28316 15487
rect 29276 15512 29328 15564
rect 29552 15555 29604 15564
rect 29552 15521 29561 15555
rect 29561 15521 29595 15555
rect 29595 15521 29604 15555
rect 29552 15512 29604 15521
rect 31668 15555 31720 15564
rect 31668 15521 31677 15555
rect 31677 15521 31711 15555
rect 31711 15521 31720 15555
rect 31668 15512 31720 15521
rect 28264 15444 28316 15453
rect 28816 15444 28868 15496
rect 30656 15444 30708 15496
rect 29368 15308 29420 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9680 15104 9732 15156
rect 13452 15104 13504 15156
rect 21548 15104 21600 15156
rect 22008 15104 22060 15156
rect 23572 15104 23624 15156
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 10232 15036 10284 15088
rect 17960 15036 18012 15088
rect 11888 14968 11940 15020
rect 12164 14968 12216 15020
rect 13176 14968 13228 15020
rect 14924 14968 14976 15020
rect 16948 14968 17000 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 18604 15036 18656 15088
rect 20352 15036 20404 15088
rect 22100 15036 22152 15088
rect 25596 15104 25648 15156
rect 25964 15104 26016 15156
rect 27712 15104 27764 15156
rect 30656 15147 30708 15156
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 17868 14900 17920 14952
rect 19524 14900 19576 14952
rect 20352 14900 20404 14952
rect 21272 14968 21324 15020
rect 21824 14968 21876 15020
rect 23480 14968 23532 15020
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 24952 15036 25004 15088
rect 25688 15036 25740 15088
rect 27896 15036 27948 15088
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 31208 15079 31260 15088
rect 24676 14968 24728 15020
rect 24860 14968 24912 15020
rect 25320 15011 25372 15020
rect 25320 14977 25343 15011
rect 25343 14977 25372 15011
rect 25320 14968 25372 14977
rect 26976 15011 27028 15020
rect 26976 14977 26985 15011
rect 26985 14977 27019 15011
rect 27019 14977 27028 15011
rect 26976 14968 27028 14977
rect 20812 14900 20864 14952
rect 15384 14832 15436 14884
rect 19432 14832 19484 14884
rect 19892 14832 19944 14884
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 22652 14900 22704 14952
rect 11520 14764 11572 14816
rect 13084 14764 13136 14816
rect 18052 14764 18104 14816
rect 21456 14832 21508 14884
rect 24124 14900 24176 14952
rect 26332 14900 26384 14952
rect 27988 14968 28040 15020
rect 31208 15045 31217 15079
rect 31217 15045 31251 15079
rect 31251 15045 31260 15079
rect 31208 15036 31260 15045
rect 28356 14968 28408 15020
rect 29276 15011 29328 15020
rect 29276 14977 29285 15011
rect 29285 14977 29319 15011
rect 29319 14977 29328 15011
rect 29276 14968 29328 14977
rect 29368 14968 29420 15020
rect 29184 14900 29236 14952
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 22652 14764 22704 14816
rect 25044 14832 25096 14884
rect 23204 14764 23256 14816
rect 23480 14764 23532 14816
rect 24400 14764 24452 14816
rect 24584 14764 24636 14816
rect 28816 14832 28868 14884
rect 29644 14764 29696 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 16120 14560 16172 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 17592 14492 17644 14544
rect 19524 14492 19576 14544
rect 22284 14560 22336 14612
rect 23572 14560 23624 14612
rect 25780 14560 25832 14612
rect 26240 14560 26292 14612
rect 28264 14560 28316 14612
rect 31208 14560 31260 14612
rect 22468 14492 22520 14544
rect 25596 14492 25648 14544
rect 25964 14492 26016 14544
rect 26884 14492 26936 14544
rect 17132 14424 17184 14476
rect 17868 14424 17920 14476
rect 11336 14331 11388 14340
rect 11336 14297 11345 14331
rect 11345 14297 11379 14331
rect 11379 14297 11388 14331
rect 11336 14288 11388 14297
rect 12900 14331 12952 14340
rect 12900 14297 12909 14331
rect 12909 14297 12943 14331
rect 12943 14297 12952 14331
rect 12900 14288 12952 14297
rect 13452 14288 13504 14340
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 14372 14356 14424 14408
rect 16212 14356 16264 14408
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 18604 14424 18656 14476
rect 19984 14467 20036 14476
rect 19984 14433 19993 14467
rect 19993 14433 20027 14467
rect 20027 14433 20036 14467
rect 19984 14424 20036 14433
rect 18420 14356 18472 14408
rect 18696 14356 18748 14408
rect 19432 14356 19484 14408
rect 20628 14356 20680 14408
rect 21548 14356 21600 14408
rect 22100 14356 22152 14408
rect 22192 14356 22244 14408
rect 22652 14399 22704 14408
rect 15292 14288 15344 14340
rect 16672 14288 16724 14340
rect 20904 14288 20956 14340
rect 15660 14220 15712 14272
rect 18144 14220 18196 14272
rect 18420 14220 18472 14272
rect 22008 14220 22060 14272
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 22744 14399 22796 14408
rect 22744 14365 22754 14399
rect 22754 14365 22788 14399
rect 22788 14365 22796 14399
rect 22744 14356 22796 14365
rect 23112 14399 23164 14408
rect 23112 14365 23126 14399
rect 23126 14365 23160 14399
rect 23160 14365 23164 14399
rect 24400 14399 24452 14408
rect 23112 14356 23164 14365
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 24676 14399 24728 14408
rect 22928 14331 22980 14340
rect 22928 14297 22937 14331
rect 22937 14297 22971 14331
rect 22971 14297 22980 14331
rect 22928 14288 22980 14297
rect 23848 14288 23900 14340
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 24768 14331 24820 14340
rect 24768 14297 24777 14331
rect 24777 14297 24811 14331
rect 24811 14297 24820 14331
rect 25044 14356 25096 14408
rect 27804 14424 27856 14476
rect 28540 14424 28592 14476
rect 27620 14399 27672 14408
rect 27620 14365 27629 14399
rect 27629 14365 27663 14399
rect 27663 14365 27672 14399
rect 29276 14424 29328 14476
rect 27620 14356 27672 14365
rect 24768 14288 24820 14297
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 24860 14220 24912 14272
rect 25688 14263 25740 14272
rect 25688 14229 25713 14263
rect 25713 14229 25740 14263
rect 27712 14288 27764 14340
rect 25688 14220 25740 14229
rect 26884 14263 26936 14272
rect 26884 14229 26893 14263
rect 26893 14229 26927 14263
rect 26927 14229 26936 14263
rect 26884 14220 26936 14229
rect 27436 14220 27488 14272
rect 28908 14399 28960 14408
rect 28908 14365 28917 14399
rect 28917 14365 28951 14399
rect 28951 14365 28960 14399
rect 28908 14356 28960 14365
rect 29644 14356 29696 14408
rect 29092 14288 29144 14340
rect 28356 14220 28408 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9772 14016 9824 14068
rect 10508 13948 10560 14000
rect 11888 14016 11940 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 11796 13948 11848 14000
rect 16396 13948 16448 14000
rect 18236 14016 18288 14068
rect 10232 13880 10284 13932
rect 11336 13880 11388 13932
rect 13268 13880 13320 13932
rect 14556 13880 14608 13932
rect 15200 13880 15252 13932
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 17868 13948 17920 14000
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 17500 13880 17552 13932
rect 17592 13880 17644 13932
rect 18696 13948 18748 14000
rect 18972 13880 19024 13932
rect 15752 13812 15804 13864
rect 17960 13812 18012 13864
rect 17132 13744 17184 13796
rect 19064 13744 19116 13796
rect 20352 14016 20404 14068
rect 20628 14016 20680 14068
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 20168 13880 20220 13932
rect 20352 13880 20404 13932
rect 20812 14016 20864 14068
rect 24308 14016 24360 14068
rect 24584 14059 24636 14068
rect 24584 14025 24593 14059
rect 24593 14025 24627 14059
rect 24627 14025 24636 14059
rect 24584 14016 24636 14025
rect 22192 13948 22244 14000
rect 21732 13880 21784 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 22836 13923 22888 13932
rect 22836 13889 22845 13923
rect 22845 13889 22879 13923
rect 22879 13889 22888 13923
rect 22836 13880 22888 13889
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 29184 14016 29236 14068
rect 26056 13991 26108 14000
rect 26056 13957 26065 13991
rect 26065 13957 26099 13991
rect 26099 13957 26108 13991
rect 26056 13948 26108 13957
rect 24860 13880 24912 13889
rect 28632 13948 28684 14000
rect 28724 13948 28776 14000
rect 27436 13923 27488 13932
rect 27436 13889 27470 13923
rect 27470 13889 27488 13923
rect 27436 13880 27488 13889
rect 29184 13923 29236 13932
rect 29184 13889 29193 13923
rect 29193 13889 29227 13923
rect 29227 13889 29236 13923
rect 29184 13880 29236 13889
rect 20536 13812 20588 13864
rect 22652 13812 22704 13864
rect 22744 13812 22796 13864
rect 22928 13812 22980 13864
rect 25688 13812 25740 13864
rect 28540 13812 28592 13864
rect 20076 13744 20128 13796
rect 22468 13744 22520 13796
rect 23020 13744 23072 13796
rect 23204 13744 23256 13796
rect 24676 13744 24728 13796
rect 24860 13744 24912 13796
rect 25136 13744 25188 13796
rect 11060 13676 11112 13728
rect 14280 13719 14332 13728
rect 14280 13685 14289 13719
rect 14289 13685 14323 13719
rect 14323 13685 14332 13719
rect 14280 13676 14332 13685
rect 17684 13676 17736 13728
rect 17868 13676 17920 13728
rect 18696 13676 18748 13728
rect 18880 13676 18932 13728
rect 19248 13676 19300 13728
rect 19616 13676 19668 13728
rect 20260 13676 20312 13728
rect 23388 13676 23440 13728
rect 25228 13676 25280 13728
rect 25320 13676 25372 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 26976 13676 27028 13728
rect 29000 13719 29052 13728
rect 29000 13685 29009 13719
rect 29009 13685 29043 13719
rect 29043 13685 29052 13719
rect 29000 13676 29052 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10968 13472 11020 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 13360 13447 13412 13456
rect 13360 13413 13369 13447
rect 13369 13413 13403 13447
rect 13403 13413 13412 13447
rect 13360 13404 13412 13413
rect 17224 13447 17276 13456
rect 17224 13413 17233 13447
rect 17233 13413 17267 13447
rect 17267 13413 17276 13447
rect 17224 13404 17276 13413
rect 17684 13404 17736 13456
rect 9036 13268 9088 13320
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 9772 13311 9824 13320
rect 9772 13277 9806 13311
rect 9806 13277 9824 13311
rect 9772 13268 9824 13277
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 11980 13268 12032 13320
rect 19432 13336 19484 13388
rect 11336 13243 11388 13252
rect 11336 13209 11345 13243
rect 11345 13209 11379 13243
rect 11379 13209 11388 13243
rect 11336 13200 11388 13209
rect 12992 13200 13044 13252
rect 13636 13268 13688 13320
rect 14004 13268 14056 13320
rect 14464 13268 14516 13320
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 15844 13268 15896 13320
rect 18144 13268 18196 13320
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 19340 13268 19392 13320
rect 19984 13472 20036 13524
rect 20996 13472 21048 13524
rect 23112 13472 23164 13524
rect 22100 13336 22152 13388
rect 21272 13268 21324 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 22928 13336 22980 13388
rect 24492 13472 24544 13524
rect 26424 13472 26476 13524
rect 24216 13404 24268 13456
rect 24124 13336 24176 13388
rect 24768 13404 24820 13456
rect 26884 13404 26936 13456
rect 24400 13311 24452 13320
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13820 13132 13872 13184
rect 14740 13175 14792 13184
rect 14740 13141 14749 13175
rect 14749 13141 14783 13175
rect 14783 13141 14792 13175
rect 14740 13132 14792 13141
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 15936 13132 15988 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 20076 13200 20128 13252
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 24952 13336 25004 13388
rect 24860 13311 24912 13320
rect 24860 13277 24874 13311
rect 24874 13277 24908 13311
rect 24908 13277 24912 13311
rect 24860 13268 24912 13277
rect 25596 13268 25648 13320
rect 29184 13472 29236 13524
rect 29092 13404 29144 13456
rect 27252 13268 27304 13320
rect 26424 13200 26476 13252
rect 20628 13132 20680 13184
rect 22468 13132 22520 13184
rect 23020 13132 23072 13184
rect 27528 13132 27580 13184
rect 27712 13200 27764 13252
rect 28816 13311 28868 13320
rect 28816 13277 28825 13311
rect 28825 13277 28859 13311
rect 28859 13277 28868 13311
rect 28816 13268 28868 13277
rect 27896 13200 27948 13252
rect 28908 13132 28960 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 10232 12971 10284 12980
rect 10232 12937 10241 12971
rect 10241 12937 10275 12971
rect 10275 12937 10284 12971
rect 10232 12928 10284 12937
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 14004 12928 14056 12980
rect 14464 12928 14516 12980
rect 14832 12971 14884 12980
rect 14832 12937 14841 12971
rect 14841 12937 14875 12971
rect 14875 12937 14884 12971
rect 14832 12928 14884 12937
rect 17040 12928 17092 12980
rect 20076 12971 20128 12980
rect 12440 12860 12492 12912
rect 14740 12860 14792 12912
rect 16948 12860 17000 12912
rect 11060 12792 11112 12844
rect 12164 12792 12216 12844
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 15752 12792 15804 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18236 12860 18288 12912
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 21088 12928 21140 12980
rect 19432 12792 19484 12844
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 20628 12792 20680 12844
rect 21272 12835 21324 12844
rect 11428 12724 11480 12776
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 18052 12724 18104 12776
rect 10968 12656 11020 12708
rect 12992 12588 13044 12640
rect 16212 12656 16264 12708
rect 20996 12724 21048 12776
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 21640 12724 21692 12776
rect 22468 12928 22520 12980
rect 22836 12860 22888 12912
rect 23480 12928 23532 12980
rect 23756 12860 23808 12912
rect 25504 12860 25556 12912
rect 25688 12903 25740 12912
rect 25688 12869 25697 12903
rect 25697 12869 25731 12903
rect 25731 12869 25740 12903
rect 25688 12860 25740 12869
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 23020 12835 23072 12844
rect 22008 12792 22060 12801
rect 23020 12801 23054 12835
rect 23054 12801 23072 12835
rect 23020 12792 23072 12801
rect 22468 12724 22520 12776
rect 24400 12792 24452 12844
rect 19340 12656 19392 12708
rect 20168 12656 20220 12708
rect 21180 12656 21232 12708
rect 24124 12699 24176 12708
rect 24124 12665 24133 12699
rect 24133 12665 24167 12699
rect 24167 12665 24176 12699
rect 24124 12656 24176 12665
rect 24676 12656 24728 12708
rect 26424 12860 26476 12912
rect 29000 12860 29052 12912
rect 26976 12835 27028 12844
rect 26976 12801 26985 12835
rect 26985 12801 27019 12835
rect 27019 12801 27028 12835
rect 26976 12792 27028 12801
rect 25228 12724 25280 12776
rect 27620 12792 27672 12844
rect 28632 12835 28684 12844
rect 28632 12801 28641 12835
rect 28641 12801 28675 12835
rect 28675 12801 28684 12835
rect 28632 12792 28684 12801
rect 24860 12656 24912 12708
rect 25044 12656 25096 12708
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 20536 12588 20588 12640
rect 23112 12588 23164 12640
rect 24216 12588 24268 12640
rect 25320 12588 25372 12640
rect 27252 12656 27304 12708
rect 26148 12588 26200 12640
rect 27896 12588 27948 12640
rect 28816 12588 28868 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 11336 12384 11388 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 14924 12384 14976 12436
rect 16028 12384 16080 12436
rect 9956 12180 10008 12232
rect 11796 12248 11848 12300
rect 13728 12248 13780 12300
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 14004 12180 14056 12232
rect 12440 12112 12492 12164
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 10600 12044 10652 12096
rect 12992 12044 13044 12096
rect 14832 12180 14884 12232
rect 15568 12180 15620 12232
rect 17500 12180 17552 12232
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 15016 12112 15068 12164
rect 16120 12112 16172 12164
rect 20628 12359 20680 12368
rect 20628 12325 20637 12359
rect 20637 12325 20671 12359
rect 20671 12325 20680 12359
rect 20628 12316 20680 12325
rect 24216 12316 24268 12368
rect 25044 12384 25096 12436
rect 27160 12316 27212 12368
rect 27620 12291 27672 12300
rect 22744 12180 22796 12232
rect 23112 12180 23164 12232
rect 23388 12180 23440 12232
rect 19984 12112 20036 12164
rect 20260 12112 20312 12164
rect 23480 12112 23532 12164
rect 16304 12044 16356 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 21180 12044 21232 12096
rect 23204 12044 23256 12096
rect 24032 12180 24084 12232
rect 24492 12180 24544 12232
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 27620 12257 27629 12291
rect 27629 12257 27663 12291
rect 27663 12257 27672 12291
rect 27620 12248 27672 12257
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 27252 12180 27304 12232
rect 28172 12180 28224 12232
rect 25964 12112 26016 12164
rect 24860 12044 24912 12096
rect 25228 12044 25280 12096
rect 25596 12044 25648 12096
rect 26700 12044 26752 12096
rect 28448 12112 28500 12164
rect 29552 12087 29604 12096
rect 29552 12053 29561 12087
rect 29561 12053 29595 12087
rect 29595 12053 29604 12087
rect 29552 12044 29604 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 11428 11840 11480 11892
rect 14188 11840 14240 11892
rect 15108 11840 15160 11892
rect 15200 11840 15252 11892
rect 17592 11840 17644 11892
rect 20260 11883 20312 11892
rect 20260 11849 20269 11883
rect 20269 11849 20303 11883
rect 20303 11849 20312 11883
rect 20260 11840 20312 11849
rect 20720 11840 20772 11892
rect 22836 11840 22888 11892
rect 24032 11840 24084 11892
rect 8944 11772 8996 11824
rect 8852 11704 8904 11756
rect 11888 11704 11940 11756
rect 12256 11704 12308 11756
rect 12992 11747 13044 11756
rect 12992 11713 13026 11747
rect 13026 11713 13044 11747
rect 12992 11704 13044 11713
rect 18052 11772 18104 11824
rect 15292 11704 15344 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 20996 11772 21048 11824
rect 6552 11636 6604 11688
rect 8484 11636 8536 11688
rect 9036 11636 9088 11688
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 10600 11636 10652 11688
rect 15660 11636 15712 11688
rect 18052 11636 18104 11688
rect 19064 11704 19116 11756
rect 20720 11704 20772 11756
rect 21180 11772 21232 11824
rect 19248 11636 19300 11688
rect 23848 11772 23900 11824
rect 25412 11840 25464 11892
rect 24492 11772 24544 11824
rect 22008 11704 22060 11756
rect 23388 11747 23440 11756
rect 23388 11713 23397 11747
rect 23397 11713 23431 11747
rect 23431 11713 23440 11747
rect 23388 11704 23440 11713
rect 21456 11636 21508 11688
rect 18512 11568 18564 11620
rect 18972 11568 19024 11620
rect 6276 11500 6328 11552
rect 9036 11500 9088 11552
rect 9588 11500 9640 11552
rect 16580 11500 16632 11552
rect 17592 11500 17644 11552
rect 17868 11500 17920 11552
rect 18696 11500 18748 11552
rect 19340 11500 19392 11552
rect 22008 11568 22060 11620
rect 22192 11500 22244 11552
rect 24860 11636 24912 11688
rect 25228 11772 25280 11824
rect 28172 11840 28224 11892
rect 28908 11840 28960 11892
rect 25872 11772 25924 11824
rect 27712 11772 27764 11824
rect 29552 11772 29604 11824
rect 25964 11704 26016 11756
rect 27528 11704 27580 11756
rect 28632 11704 28684 11756
rect 28264 11636 28316 11688
rect 24584 11568 24636 11620
rect 24952 11500 25004 11552
rect 25044 11500 25096 11552
rect 26516 11500 26568 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 8852 11296 8904 11348
rect 9036 11296 9088 11348
rect 7656 11228 7708 11280
rect 12624 11228 12676 11280
rect 15476 11296 15528 11348
rect 16672 11296 16724 11348
rect 16856 11296 16908 11348
rect 17040 11296 17092 11348
rect 17316 11296 17368 11348
rect 17500 11296 17552 11348
rect 20812 11296 20864 11348
rect 20904 11296 20956 11348
rect 23204 11296 23256 11348
rect 23480 11296 23532 11348
rect 24860 11296 24912 11348
rect 25872 11296 25924 11348
rect 28448 11339 28500 11348
rect 4896 11092 4948 11144
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 8392 11092 8444 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9404 11092 9456 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 13728 11092 13780 11144
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 16028 11092 16080 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 16580 11135 16632 11144
rect 16580 11101 16613 11135
rect 16613 11101 16632 11135
rect 16580 11092 16632 11101
rect 16856 11092 16908 11144
rect 17868 11228 17920 11280
rect 20628 11271 20680 11280
rect 20628 11237 20637 11271
rect 20637 11237 20671 11271
rect 20671 11237 20680 11271
rect 20628 11228 20680 11237
rect 21180 11228 21232 11280
rect 21548 11228 21600 11280
rect 26240 11228 26292 11280
rect 21732 11203 21784 11212
rect 6644 11024 6696 11076
rect 10048 11067 10100 11076
rect 10048 11033 10082 11067
rect 10082 11033 10100 11067
rect 10048 11024 10100 11033
rect 10968 11024 11020 11076
rect 15016 11024 15068 11076
rect 10692 10956 10744 11008
rect 16120 11024 16172 11076
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17868 11092 17920 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18512 11092 18564 11144
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 22284 11160 22336 11212
rect 20996 11092 21048 11144
rect 21456 11092 21508 11144
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 24676 11160 24728 11212
rect 21548 11092 21600 11101
rect 23112 11092 23164 11144
rect 23388 11092 23440 11144
rect 15660 10956 15712 11008
rect 16856 10956 16908 11008
rect 17040 10956 17092 11008
rect 21088 11024 21140 11076
rect 21824 11024 21876 11076
rect 22100 11024 22152 11076
rect 23848 11092 23900 11144
rect 25596 11160 25648 11212
rect 25780 11160 25832 11212
rect 26424 11160 26476 11212
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 24584 11024 24636 11033
rect 25872 11135 25924 11144
rect 25872 11101 25886 11135
rect 25886 11101 25920 11135
rect 25920 11101 25924 11135
rect 26516 11135 26568 11144
rect 25872 11092 25924 11101
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 28448 11305 28457 11339
rect 28457 11305 28491 11339
rect 28491 11305 28500 11339
rect 28448 11296 28500 11305
rect 29092 11296 29144 11348
rect 31484 11339 31536 11348
rect 31484 11305 31493 11339
rect 31493 11305 31527 11339
rect 31527 11305 31536 11339
rect 31484 11296 31536 11305
rect 27160 11271 27212 11280
rect 27160 11237 27169 11271
rect 27169 11237 27203 11271
rect 27203 11237 27212 11271
rect 27160 11228 27212 11237
rect 27344 11228 27396 11280
rect 26884 11160 26936 11212
rect 27712 11092 27764 11144
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 28724 11092 28776 11144
rect 29552 11092 29604 11144
rect 26240 11024 26292 11076
rect 26332 11024 26384 11076
rect 26424 11024 26476 11076
rect 23204 10956 23256 11008
rect 28080 11024 28132 11076
rect 29828 11092 29880 11144
rect 28908 10956 28960 11008
rect 29552 10999 29604 11008
rect 29552 10965 29561 10999
rect 29561 10965 29595 10999
rect 29595 10965 29604 10999
rect 29552 10956 29604 10965
rect 30840 10999 30892 11008
rect 30840 10965 30849 10999
rect 30849 10965 30883 10999
rect 30883 10965 30892 10999
rect 30840 10956 30892 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 6644 10752 6696 10804
rect 9128 10752 9180 10804
rect 9956 10752 10008 10804
rect 11796 10752 11848 10804
rect 14004 10752 14056 10804
rect 18236 10752 18288 10804
rect 20444 10752 20496 10804
rect 7012 10616 7064 10668
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 1584 10480 1636 10532
rect 6736 10412 6788 10464
rect 8392 10412 8444 10464
rect 15016 10684 15068 10736
rect 21916 10684 21968 10736
rect 11704 10659 11756 10668
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 15108 10659 15160 10668
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 11060 10480 11112 10532
rect 12900 10548 12952 10600
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15568 10616 15620 10668
rect 17040 10616 17092 10668
rect 18144 10616 18196 10668
rect 16580 10548 16632 10600
rect 11152 10412 11204 10464
rect 17868 10548 17920 10600
rect 19248 10616 19300 10668
rect 20076 10616 20128 10668
rect 20904 10616 20956 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 21180 10616 21232 10668
rect 19984 10548 20036 10600
rect 20720 10548 20772 10600
rect 21548 10616 21600 10668
rect 22008 10616 22060 10668
rect 23664 10727 23716 10736
rect 23664 10693 23673 10727
rect 23673 10693 23707 10727
rect 23707 10693 23716 10727
rect 23664 10684 23716 10693
rect 21456 10548 21508 10600
rect 23756 10659 23808 10668
rect 23204 10548 23256 10600
rect 23756 10625 23765 10659
rect 23765 10625 23799 10659
rect 23799 10625 23808 10659
rect 23756 10616 23808 10625
rect 24860 10659 24912 10668
rect 24860 10625 24869 10659
rect 24869 10625 24903 10659
rect 24903 10625 24912 10659
rect 24860 10616 24912 10625
rect 25780 10616 25832 10668
rect 24492 10548 24544 10600
rect 25228 10548 25280 10600
rect 28908 10752 28960 10804
rect 27620 10616 27672 10668
rect 29552 10616 29604 10668
rect 30472 10616 30524 10668
rect 31576 10659 31628 10668
rect 20168 10480 20220 10532
rect 20996 10480 21048 10532
rect 22100 10480 22152 10532
rect 22744 10480 22796 10532
rect 23664 10480 23716 10532
rect 27528 10480 27580 10532
rect 17408 10412 17460 10464
rect 19340 10412 19392 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 21088 10412 21140 10464
rect 23848 10412 23900 10464
rect 27068 10412 27120 10464
rect 28724 10548 28776 10600
rect 31576 10625 31585 10659
rect 31585 10625 31619 10659
rect 31619 10625 31628 10659
rect 31576 10616 31628 10625
rect 31300 10480 31352 10532
rect 30840 10412 30892 10464
rect 31024 10412 31076 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6552 10208 6604 10260
rect 7012 10208 7064 10260
rect 9772 10208 9824 10260
rect 11244 10208 11296 10260
rect 11704 10208 11756 10260
rect 12072 10208 12124 10260
rect 13912 10208 13964 10260
rect 15108 10208 15160 10260
rect 16948 10208 17000 10260
rect 18420 10208 18472 10260
rect 5264 10140 5316 10192
rect 7104 10072 7156 10124
rect 11060 10072 11112 10124
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 6644 10004 6696 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8116 10004 8168 10056
rect 6920 9936 6972 9988
rect 9496 9936 9548 9988
rect 10692 10004 10744 10056
rect 11244 10072 11296 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 15568 10115 15620 10124
rect 14096 10072 14148 10081
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 16120 10072 16172 10124
rect 19064 10140 19116 10192
rect 19524 10183 19576 10192
rect 19524 10149 19533 10183
rect 19533 10149 19567 10183
rect 19567 10149 19576 10183
rect 19524 10140 19576 10149
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 21548 10208 21600 10260
rect 19984 10140 20036 10192
rect 23756 10208 23808 10260
rect 26240 10251 26292 10260
rect 26240 10217 26249 10251
rect 26249 10217 26283 10251
rect 26283 10217 26292 10251
rect 26240 10208 26292 10217
rect 26424 10208 26476 10260
rect 27344 10140 27396 10192
rect 17868 10072 17920 10124
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 12072 10004 12124 10056
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 11060 9936 11112 9988
rect 11428 9936 11480 9988
rect 11612 9936 11664 9988
rect 12808 9936 12860 9988
rect 13912 10004 13964 10056
rect 15384 10004 15436 10056
rect 16488 10004 16540 10056
rect 19340 10072 19392 10124
rect 20076 10072 20128 10124
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 16856 9936 16908 9988
rect 18420 9936 18472 9988
rect 20996 10004 21048 10056
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 23480 10004 23532 10056
rect 24492 10004 24544 10056
rect 20444 9936 20496 9988
rect 20720 9979 20772 9988
rect 20720 9945 20729 9979
rect 20729 9945 20763 9979
rect 20763 9945 20772 9979
rect 20720 9936 20772 9945
rect 21088 9936 21140 9988
rect 23848 9936 23900 9988
rect 26240 10004 26292 10056
rect 27252 10072 27304 10124
rect 28724 10072 28776 10124
rect 27712 10004 27764 10056
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 29000 10004 29052 10013
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 30012 10072 30064 10124
rect 29828 10004 29880 10056
rect 31392 10004 31444 10056
rect 27896 9936 27948 9988
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 28172 9936 28224 9945
rect 30932 9936 30984 9988
rect 6000 9868 6052 9920
rect 9036 9868 9088 9920
rect 12072 9868 12124 9920
rect 15108 9868 15160 9920
rect 18880 9868 18932 9920
rect 19340 9868 19392 9920
rect 20260 9868 20312 9920
rect 26700 9868 26752 9920
rect 30196 9911 30248 9920
rect 30196 9877 30205 9911
rect 30205 9877 30239 9911
rect 30239 9877 30248 9911
rect 30196 9868 30248 9877
rect 30288 9868 30340 9920
rect 31484 9911 31536 9920
rect 31484 9877 31493 9911
rect 31493 9877 31527 9911
rect 31527 9877 31536 9911
rect 31484 9868 31536 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4896 9596 4948 9648
rect 7748 9664 7800 9716
rect 9496 9664 9548 9716
rect 5908 9596 5960 9648
rect 4988 9528 5040 9580
rect 5356 9528 5408 9580
rect 8576 9596 8628 9648
rect 9312 9596 9364 9648
rect 10784 9639 10836 9648
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 6276 9528 6328 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6644 9528 6696 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 6184 9460 6236 9512
rect 7748 9460 7800 9512
rect 8576 9460 8628 9512
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 11060 9528 11112 9580
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 12348 9596 12400 9648
rect 13728 9664 13780 9716
rect 16580 9664 16632 9716
rect 16672 9664 16724 9716
rect 16856 9664 16908 9716
rect 14280 9596 14332 9648
rect 12808 9528 12860 9580
rect 15200 9596 15252 9648
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 12256 9503 12308 9512
rect 6460 9392 6512 9444
rect 9128 9392 9180 9444
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 13360 9460 13412 9512
rect 15200 9460 15252 9512
rect 15660 9528 15712 9580
rect 16488 9460 16540 9512
rect 10968 9435 11020 9444
rect 10968 9401 10977 9435
rect 10977 9401 11011 9435
rect 11011 9401 11020 9435
rect 10968 9392 11020 9401
rect 5540 9324 5592 9376
rect 9036 9324 9088 9376
rect 14464 9392 14516 9444
rect 19524 9596 19576 9648
rect 21916 9664 21968 9716
rect 22376 9664 22428 9716
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17960 9528 18012 9580
rect 18236 9528 18288 9580
rect 17500 9460 17552 9512
rect 18604 9528 18656 9580
rect 19340 9528 19392 9580
rect 20444 9528 20496 9580
rect 21088 9596 21140 9648
rect 21180 9596 21232 9648
rect 22284 9596 22336 9648
rect 19064 9460 19116 9512
rect 21732 9528 21784 9580
rect 23756 9596 23808 9648
rect 24676 9528 24728 9580
rect 24952 9571 25004 9580
rect 25228 9664 25280 9716
rect 27896 9664 27948 9716
rect 25596 9596 25648 9648
rect 25688 9596 25740 9648
rect 26332 9596 26384 9648
rect 26608 9596 26660 9648
rect 26884 9596 26936 9648
rect 27068 9596 27120 9648
rect 30104 9596 30156 9648
rect 24952 9537 24968 9571
rect 24968 9537 25002 9571
rect 25002 9537 25004 9571
rect 24952 9528 25004 9537
rect 25417 9537 25426 9564
rect 25426 9537 25460 9564
rect 25460 9537 25469 9564
rect 25417 9512 25469 9537
rect 26792 9528 26844 9580
rect 27344 9571 27396 9580
rect 27344 9537 27353 9571
rect 27353 9537 27387 9571
rect 27387 9537 27396 9571
rect 27344 9528 27396 9537
rect 21088 9460 21140 9512
rect 22284 9503 22336 9512
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 20904 9392 20956 9444
rect 23664 9460 23716 9512
rect 24860 9460 24912 9512
rect 30380 9528 30432 9580
rect 30748 9596 30800 9648
rect 30564 9528 30616 9580
rect 25228 9392 25280 9444
rect 13728 9324 13780 9376
rect 14924 9324 14976 9376
rect 17224 9324 17276 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 17960 9324 18012 9376
rect 18880 9324 18932 9376
rect 22100 9324 22152 9376
rect 22192 9367 22244 9376
rect 22192 9333 22201 9367
rect 22201 9333 22235 9367
rect 22235 9333 22244 9367
rect 22192 9324 22244 9333
rect 23020 9324 23072 9376
rect 25780 9392 25832 9444
rect 26056 9392 26108 9444
rect 27620 9460 27672 9512
rect 28448 9460 28500 9512
rect 29644 9460 29696 9512
rect 31944 9528 31996 9580
rect 33600 9571 33652 9580
rect 33600 9537 33609 9571
rect 33609 9537 33643 9571
rect 33643 9537 33652 9571
rect 33600 9528 33652 9537
rect 26792 9324 26844 9376
rect 28172 9392 28224 9444
rect 27620 9324 27672 9376
rect 31484 9392 31536 9444
rect 30840 9324 30892 9376
rect 31116 9367 31168 9376
rect 31116 9333 31125 9367
rect 31125 9333 31159 9367
rect 31159 9333 31168 9367
rect 31116 9324 31168 9333
rect 31760 9324 31812 9376
rect 32496 9324 32548 9376
rect 33508 9324 33560 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3976 9120 4028 9172
rect 7288 9120 7340 9172
rect 7748 9120 7800 9172
rect 13452 9120 13504 9172
rect 13912 9120 13964 9172
rect 14280 9120 14332 9172
rect 18512 9120 18564 9172
rect 18604 9120 18656 9172
rect 19340 9163 19392 9172
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 19800 9120 19852 9172
rect 20076 9120 20128 9172
rect 20996 9120 21048 9172
rect 21364 9120 21416 9172
rect 22284 9120 22336 9172
rect 22376 9120 22428 9172
rect 3884 8916 3936 8968
rect 4160 8848 4212 8900
rect 4712 8848 4764 8900
rect 3424 8780 3476 8832
rect 11980 9052 12032 9104
rect 12348 9052 12400 9104
rect 12808 9052 12860 9104
rect 13176 9052 13228 9104
rect 6276 8916 6328 8968
rect 5172 8848 5224 8900
rect 5724 8780 5776 8832
rect 6092 8780 6144 8832
rect 6552 8848 6604 8900
rect 6736 8984 6788 9036
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 9404 8984 9456 9036
rect 6828 8916 6880 8925
rect 7748 8916 7800 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 9956 8916 10008 8968
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10324 8959 10376 8968
rect 10048 8916 10100 8925
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 11060 8916 11112 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11796 8916 11848 8968
rect 12256 8984 12308 9036
rect 12440 8916 12492 8968
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 8760 8848 8812 8900
rect 8024 8780 8076 8832
rect 10876 8780 10928 8832
rect 13636 8916 13688 8968
rect 16948 8916 17000 8968
rect 17040 8916 17092 8968
rect 17684 8916 17736 8968
rect 18328 8984 18380 9036
rect 21824 9052 21876 9104
rect 22652 9120 22704 9172
rect 23020 9120 23072 9172
rect 25596 9120 25648 9172
rect 29828 9120 29880 9172
rect 30380 9120 30432 9172
rect 18880 8984 18932 9036
rect 19800 8984 19852 9036
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 19248 8916 19300 8968
rect 19432 8916 19484 8968
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 20444 8984 20496 9036
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 11980 8780 12032 8832
rect 13176 8891 13228 8900
rect 13176 8857 13185 8891
rect 13185 8857 13219 8891
rect 13219 8857 13228 8891
rect 13176 8848 13228 8857
rect 12900 8780 12952 8832
rect 12992 8780 13044 8832
rect 13728 8780 13780 8832
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 15660 8780 15712 8789
rect 17500 8848 17552 8900
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 19064 8848 19116 8900
rect 20996 8916 21048 8968
rect 21180 8916 21232 8968
rect 22192 8916 22244 8968
rect 20812 8848 20864 8900
rect 21732 8848 21784 8900
rect 21916 8848 21968 8900
rect 23020 8916 23072 8968
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 22744 8848 22796 8900
rect 24492 9027 24544 9036
rect 24492 8993 24501 9027
rect 24501 8993 24535 9027
rect 24535 8993 24544 9027
rect 24492 8984 24544 8993
rect 31116 9052 31168 9104
rect 32220 9052 32272 9104
rect 27436 8984 27488 9036
rect 28908 9027 28960 9036
rect 28908 8993 28917 9027
rect 28917 8993 28951 9027
rect 28951 8993 28960 9027
rect 28908 8984 28960 8993
rect 29000 8984 29052 9036
rect 29184 8984 29236 9036
rect 26884 8916 26936 8968
rect 27252 8916 27304 8968
rect 27528 8916 27580 8968
rect 27068 8891 27120 8900
rect 27068 8857 27077 8891
rect 27077 8857 27111 8891
rect 27111 8857 27120 8891
rect 27068 8848 27120 8857
rect 28356 8916 28408 8968
rect 29368 8916 29420 8968
rect 29920 8916 29972 8968
rect 30380 8959 30432 8968
rect 30380 8925 30389 8959
rect 30389 8925 30423 8959
rect 30423 8925 30432 8959
rect 30380 8916 30432 8925
rect 30932 8916 30984 8968
rect 31116 8916 31168 8968
rect 32312 8959 32364 8968
rect 32312 8925 32321 8959
rect 32321 8925 32355 8959
rect 32355 8925 32364 8959
rect 32312 8916 32364 8925
rect 32956 8959 33008 8968
rect 32956 8925 32965 8959
rect 32965 8925 32999 8959
rect 32999 8925 33008 8959
rect 32956 8916 33008 8925
rect 33876 8916 33928 8968
rect 29000 8848 29052 8900
rect 18696 8780 18748 8832
rect 20260 8780 20312 8832
rect 20904 8780 20956 8832
rect 21180 8780 21232 8832
rect 21824 8780 21876 8832
rect 24400 8780 24452 8832
rect 26240 8780 26292 8832
rect 27344 8823 27396 8832
rect 27344 8789 27353 8823
rect 27353 8789 27387 8823
rect 27387 8789 27396 8823
rect 27344 8780 27396 8789
rect 28172 8780 28224 8832
rect 29460 8780 29512 8832
rect 29644 8823 29696 8832
rect 29644 8789 29653 8823
rect 29653 8789 29687 8823
rect 29687 8789 29696 8823
rect 29644 8780 29696 8789
rect 29828 8780 29880 8832
rect 32128 8823 32180 8832
rect 32128 8789 32137 8823
rect 32137 8789 32171 8823
rect 32171 8789 32180 8823
rect 32128 8780 32180 8789
rect 32772 8823 32824 8832
rect 32772 8789 32781 8823
rect 32781 8789 32815 8823
rect 32815 8789 32824 8823
rect 32772 8780 32824 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3240 8576 3292 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 5264 8508 5316 8560
rect 6644 8576 6696 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 7012 8576 7064 8628
rect 6276 8508 6328 8560
rect 6552 8551 6604 8560
rect 6552 8517 6561 8551
rect 6561 8517 6595 8551
rect 6595 8517 6604 8551
rect 6552 8508 6604 8517
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5632 8440 5684 8492
rect 6092 8440 6144 8492
rect 6644 8483 6696 8492
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 6828 8440 6880 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8392 8508 8444 8560
rect 9956 8576 10008 8628
rect 11060 8576 11112 8628
rect 12624 8576 12676 8628
rect 18052 8576 18104 8628
rect 19432 8619 19484 8628
rect 8116 8440 8168 8492
rect 5540 8372 5592 8381
rect 3792 8304 3844 8356
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 5448 8304 5500 8356
rect 7380 8347 7432 8356
rect 2964 8236 3016 8288
rect 5356 8236 5408 8288
rect 7380 8313 7389 8347
rect 7389 8313 7423 8347
rect 7423 8313 7432 8347
rect 7380 8304 7432 8313
rect 7840 8304 7892 8356
rect 6920 8236 6972 8288
rect 7932 8236 7984 8288
rect 9036 8236 9088 8288
rect 9312 8236 9364 8288
rect 11244 8508 11296 8560
rect 11704 8551 11756 8560
rect 11704 8517 11713 8551
rect 11713 8517 11747 8551
rect 11747 8517 11756 8551
rect 11704 8508 11756 8517
rect 12716 8508 12768 8560
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10324 8440 10376 8492
rect 11152 8440 11204 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 11612 8440 11664 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12808 8483 12860 8492
rect 11060 8372 11112 8424
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13636 8508 13688 8560
rect 17408 8508 17460 8560
rect 17592 8508 17644 8560
rect 18512 8508 18564 8560
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 20260 8508 20312 8560
rect 13544 8440 13596 8492
rect 15200 8440 15252 8492
rect 16212 8440 16264 8492
rect 16948 8440 17000 8492
rect 19064 8483 19116 8492
rect 9496 8304 9548 8356
rect 12532 8304 12584 8356
rect 14004 8372 14056 8424
rect 14280 8372 14332 8424
rect 15384 8372 15436 8424
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 19892 8440 19944 8492
rect 21824 8576 21876 8628
rect 23112 8576 23164 8628
rect 25044 8619 25096 8628
rect 25044 8585 25053 8619
rect 25053 8585 25087 8619
rect 25087 8585 25096 8619
rect 25044 8576 25096 8585
rect 28540 8576 28592 8628
rect 30472 8619 30524 8628
rect 30472 8585 30481 8619
rect 30481 8585 30515 8619
rect 30515 8585 30524 8619
rect 30472 8576 30524 8585
rect 30656 8576 30708 8628
rect 21732 8508 21784 8560
rect 20904 8483 20956 8492
rect 20904 8449 20913 8483
rect 20913 8449 20947 8483
rect 20947 8449 20956 8483
rect 20904 8440 20956 8449
rect 23020 8508 23072 8560
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 25872 8508 25924 8560
rect 26056 8508 26108 8560
rect 20628 8372 20680 8424
rect 12900 8304 12952 8356
rect 14096 8304 14148 8356
rect 16672 8304 16724 8356
rect 11060 8236 11112 8288
rect 12440 8236 12492 8288
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 14464 8236 14516 8288
rect 18236 8236 18288 8288
rect 18880 8304 18932 8356
rect 19984 8304 20036 8356
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 23480 8440 23532 8492
rect 24124 8440 24176 8492
rect 26240 8483 26292 8492
rect 26240 8449 26249 8483
rect 26249 8449 26283 8483
rect 26283 8449 26292 8483
rect 26240 8440 26292 8449
rect 27160 8483 27212 8492
rect 23020 8372 23072 8424
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 27896 8508 27948 8560
rect 28908 8508 28960 8560
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 30196 8440 30248 8492
rect 22652 8304 22704 8356
rect 27068 8372 27120 8424
rect 27528 8372 27580 8424
rect 24216 8347 24268 8356
rect 20444 8236 20496 8288
rect 20720 8236 20772 8288
rect 21272 8236 21324 8288
rect 21364 8236 21416 8288
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 21824 8236 21876 8245
rect 23020 8236 23072 8288
rect 24216 8313 24225 8347
rect 24225 8313 24259 8347
rect 24259 8313 24268 8347
rect 24216 8304 24268 8313
rect 24952 8304 25004 8356
rect 28080 8304 28132 8356
rect 29828 8372 29880 8424
rect 26056 8236 26108 8288
rect 28172 8236 28224 8288
rect 28816 8236 28868 8288
rect 29736 8304 29788 8356
rect 30656 8440 30708 8492
rect 33784 8576 33836 8628
rect 33232 8440 33284 8492
rect 33416 8440 33468 8492
rect 35348 8440 35400 8492
rect 30196 8236 30248 8288
rect 31852 8304 31904 8356
rect 34060 8304 34112 8356
rect 34520 8304 34572 8356
rect 32864 8236 32916 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4896 8032 4948 8084
rect 6000 8032 6052 8084
rect 6368 8032 6420 8084
rect 7840 8032 7892 8084
rect 7932 8032 7984 8084
rect 9772 8032 9824 8084
rect 11152 8032 11204 8084
rect 1308 7828 1360 7880
rect 2872 7828 2924 7880
rect 3516 7828 3568 7880
rect 4528 7828 4580 7880
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 6000 7896 6052 7948
rect 1952 7692 2004 7744
rect 3332 7692 3384 7744
rect 5080 7692 5132 7744
rect 5724 7828 5776 7880
rect 5356 7760 5408 7812
rect 6828 7828 6880 7880
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 6552 7760 6604 7812
rect 8944 7828 8996 7880
rect 8392 7760 8444 7812
rect 6920 7692 6972 7744
rect 7288 7692 7340 7744
rect 9128 7692 9180 7744
rect 16212 8032 16264 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 20168 8032 20220 8084
rect 21364 8032 21416 8084
rect 23480 8075 23532 8084
rect 12532 7828 12584 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14464 7828 14516 7880
rect 15384 7964 15436 8016
rect 16028 7964 16080 8016
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 24584 8032 24636 8084
rect 27252 8032 27304 8084
rect 27528 8032 27580 8084
rect 29184 8032 29236 8084
rect 24124 7964 24176 8016
rect 25136 7964 25188 8016
rect 28632 7964 28684 8016
rect 31116 8032 31168 8084
rect 33048 8032 33100 8084
rect 15292 7896 15344 7948
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15936 7828 15988 7880
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 21824 7896 21876 7948
rect 23664 7896 23716 7948
rect 23940 7896 23992 7948
rect 17592 7828 17644 7880
rect 17960 7871 18012 7880
rect 10968 7692 11020 7744
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11520 7692 11572 7744
rect 11888 7692 11940 7744
rect 16856 7803 16908 7812
rect 16856 7769 16865 7803
rect 16865 7769 16899 7803
rect 16899 7769 16908 7803
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 16856 7760 16908 7769
rect 17868 7760 17920 7812
rect 12900 7692 12952 7744
rect 14464 7692 14516 7744
rect 15568 7692 15620 7744
rect 17040 7735 17092 7744
rect 17040 7701 17049 7735
rect 17049 7701 17083 7735
rect 17083 7701 17092 7735
rect 17040 7692 17092 7701
rect 19340 7828 19392 7880
rect 19892 7828 19944 7880
rect 20076 7828 20128 7880
rect 20628 7828 20680 7880
rect 21272 7828 21324 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 19064 7760 19116 7812
rect 20260 7760 20312 7812
rect 20812 7760 20864 7812
rect 21640 7760 21692 7812
rect 22008 7760 22060 7812
rect 24216 7828 24268 7880
rect 27436 7828 27488 7880
rect 28540 7896 28592 7948
rect 29184 7896 29236 7948
rect 24676 7760 24728 7812
rect 26240 7760 26292 7812
rect 26424 7760 26476 7812
rect 27068 7760 27120 7812
rect 21180 7692 21232 7744
rect 22836 7692 22888 7744
rect 26516 7692 26568 7744
rect 27528 7692 27580 7744
rect 29000 7828 29052 7880
rect 32128 7964 32180 8016
rect 33140 7964 33192 8016
rect 28172 7760 28224 7812
rect 30656 7760 30708 7812
rect 28540 7692 28592 7744
rect 28908 7735 28960 7744
rect 28908 7701 28917 7735
rect 28917 7701 28951 7735
rect 28951 7701 28960 7735
rect 28908 7692 28960 7701
rect 29552 7692 29604 7744
rect 32036 7760 32088 7812
rect 33324 7828 33376 7880
rect 33232 7760 33284 7812
rect 34796 7828 34848 7880
rect 36084 7896 36136 7948
rect 35716 7828 35768 7880
rect 36452 7871 36504 7880
rect 36452 7837 36461 7871
rect 36461 7837 36495 7871
rect 36495 7837 36504 7871
rect 36452 7828 36504 7837
rect 36636 7828 36688 7880
rect 38016 7871 38068 7880
rect 38016 7837 38025 7871
rect 38025 7837 38059 7871
rect 38059 7837 38068 7871
rect 38016 7828 38068 7837
rect 32128 7692 32180 7744
rect 33692 7692 33744 7744
rect 34704 7735 34756 7744
rect 34704 7701 34713 7735
rect 34713 7701 34747 7735
rect 34747 7701 34756 7735
rect 34704 7692 34756 7701
rect 35440 7692 35492 7744
rect 35624 7735 35676 7744
rect 35624 7701 35633 7735
rect 35633 7701 35667 7735
rect 35667 7701 35676 7735
rect 35624 7692 35676 7701
rect 36268 7735 36320 7744
rect 36268 7701 36277 7735
rect 36277 7701 36311 7735
rect 36311 7701 36320 7735
rect 36268 7692 36320 7701
rect 37648 7692 37700 7744
rect 37832 7735 37884 7744
rect 37832 7701 37841 7735
rect 37841 7701 37875 7735
rect 37875 7701 37884 7735
rect 37832 7692 37884 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 6828 7488 6880 7540
rect 10232 7488 10284 7540
rect 940 7352 992 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 4436 7352 4488 7404
rect 3976 7284 4028 7336
rect 5356 7352 5408 7404
rect 6920 7420 6972 7472
rect 7840 7420 7892 7472
rect 11612 7488 11664 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 14280 7488 14332 7540
rect 14556 7488 14608 7540
rect 14740 7488 14792 7540
rect 15200 7531 15252 7540
rect 15200 7497 15209 7531
rect 15209 7497 15243 7531
rect 15243 7497 15252 7531
rect 15200 7488 15252 7497
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 12072 7420 12124 7472
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 7012 7352 7064 7404
rect 8484 7352 8536 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9772 7352 9824 7404
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 11060 7352 11112 7404
rect 11152 7352 11204 7404
rect 6828 7284 6880 7336
rect 6920 7284 6972 7336
rect 5172 7216 5224 7268
rect 5540 7216 5592 7268
rect 1768 7148 1820 7200
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4896 7148 4948 7200
rect 6368 7148 6420 7200
rect 8116 7148 8168 7200
rect 10048 7284 10100 7336
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 12256 7352 12308 7404
rect 12164 7284 12216 7336
rect 8300 7216 8352 7268
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9312 7148 9364 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 10232 7216 10284 7268
rect 14004 7352 14056 7404
rect 15660 7420 15712 7472
rect 16580 7420 16632 7472
rect 17592 7420 17644 7472
rect 18420 7420 18472 7472
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 14372 7284 14424 7336
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 15200 7352 15252 7404
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 17224 7352 17276 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 22100 7420 22152 7472
rect 22376 7420 22428 7472
rect 20536 7352 20588 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23020 7488 23072 7540
rect 24676 7488 24728 7540
rect 28632 7488 28684 7540
rect 24584 7420 24636 7472
rect 26884 7420 26936 7472
rect 27620 7463 27672 7472
rect 23940 7352 23992 7404
rect 24032 7352 24084 7404
rect 24768 7395 24820 7404
rect 24768 7361 24777 7395
rect 24777 7361 24811 7395
rect 24811 7361 24820 7395
rect 24768 7352 24820 7361
rect 25596 7352 25648 7404
rect 26148 7352 26200 7404
rect 26424 7395 26476 7404
rect 26424 7361 26433 7395
rect 26433 7361 26467 7395
rect 26467 7361 26476 7395
rect 26424 7352 26476 7361
rect 26516 7352 26568 7404
rect 27620 7429 27629 7463
rect 27629 7429 27663 7463
rect 27663 7429 27672 7463
rect 27620 7420 27672 7429
rect 28908 7420 28960 7472
rect 30288 7420 30340 7472
rect 28172 7352 28224 7404
rect 29184 7395 29236 7404
rect 12072 7148 12124 7200
rect 13268 7148 13320 7200
rect 14832 7216 14884 7268
rect 15108 7216 15160 7268
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 14188 7148 14240 7200
rect 29184 7361 29193 7395
rect 29193 7361 29227 7395
rect 29227 7361 29236 7395
rect 29184 7352 29236 7361
rect 31116 7420 31168 7472
rect 32312 7488 32364 7540
rect 32772 7420 32824 7472
rect 34704 7420 34756 7472
rect 36084 7420 36136 7472
rect 16488 7148 16540 7200
rect 19892 7216 19944 7268
rect 22284 7216 22336 7268
rect 23388 7216 23440 7268
rect 18604 7191 18656 7200
rect 18604 7157 18613 7191
rect 18613 7157 18647 7191
rect 18647 7157 18656 7191
rect 18604 7148 18656 7157
rect 19340 7148 19392 7200
rect 22836 7148 22888 7200
rect 24308 7148 24360 7200
rect 24400 7148 24452 7200
rect 25136 7216 25188 7268
rect 25504 7191 25556 7200
rect 25504 7157 25513 7191
rect 25513 7157 25547 7191
rect 25547 7157 25556 7191
rect 25504 7148 25556 7157
rect 28356 7216 28408 7268
rect 29552 7148 29604 7200
rect 29828 7148 29880 7200
rect 31208 7191 31260 7200
rect 31208 7157 31217 7191
rect 31217 7157 31251 7191
rect 31251 7157 31260 7191
rect 31208 7148 31260 7157
rect 33600 7352 33652 7404
rect 34796 7352 34848 7404
rect 36176 7395 36228 7404
rect 36176 7361 36185 7395
rect 36185 7361 36219 7395
rect 36219 7361 36228 7395
rect 36176 7352 36228 7361
rect 36820 7352 36872 7404
rect 36912 7352 36964 7404
rect 38108 7395 38160 7404
rect 38108 7361 38117 7395
rect 38117 7361 38151 7395
rect 38151 7361 38160 7395
rect 38108 7352 38160 7361
rect 31944 7284 31996 7336
rect 33968 7327 34020 7336
rect 33968 7293 33977 7327
rect 33977 7293 34011 7327
rect 34011 7293 34020 7327
rect 33968 7284 34020 7293
rect 36728 7216 36780 7268
rect 32128 7148 32180 7200
rect 32404 7148 32456 7200
rect 35440 7148 35492 7200
rect 35808 7191 35860 7200
rect 35808 7157 35817 7191
rect 35817 7157 35851 7191
rect 35851 7157 35860 7191
rect 35808 7148 35860 7157
rect 37280 7191 37332 7200
rect 37280 7157 37289 7191
rect 37289 7157 37323 7191
rect 37323 7157 37332 7191
rect 37280 7148 37332 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2964 6987 3016 6996
rect 2964 6953 2973 6987
rect 2973 6953 3007 6987
rect 3007 6953 3016 6987
rect 2964 6944 3016 6953
rect 3056 6944 3108 6996
rect 4528 6876 4580 6928
rect 4712 6919 4764 6928
rect 4712 6885 4721 6919
rect 4721 6885 4755 6919
rect 4755 6885 4764 6919
rect 7104 6944 7156 6996
rect 8852 6944 8904 6996
rect 9680 6944 9732 6996
rect 10600 6944 10652 6996
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 12348 6987 12400 6996
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 12440 6944 12492 6996
rect 13176 6944 13228 6996
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 15936 6944 15988 6996
rect 4712 6876 4764 6885
rect 13452 6876 13504 6928
rect 13728 6876 13780 6928
rect 3884 6808 3936 6860
rect 5448 6808 5500 6860
rect 7196 6808 7248 6860
rect 9680 6808 9732 6860
rect 9956 6808 10008 6860
rect 10692 6808 10744 6860
rect 12624 6808 12676 6860
rect 2412 6740 2464 6792
rect 2780 6740 2832 6792
rect 3240 6740 3292 6792
rect 4804 6740 4856 6792
rect 5540 6672 5592 6724
rect 5908 6672 5960 6724
rect 6552 6672 6604 6724
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 9312 6740 9364 6792
rect 9588 6740 9640 6792
rect 11244 6740 11296 6792
rect 12900 6740 12952 6792
rect 13912 6808 13964 6860
rect 19432 6944 19484 6996
rect 22652 6944 22704 6996
rect 27896 6944 27948 6996
rect 31576 6944 31628 6996
rect 13084 6740 13136 6792
rect 13636 6740 13688 6792
rect 7288 6672 7340 6724
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 4896 6604 4948 6656
rect 4988 6604 5040 6656
rect 6828 6604 6880 6656
rect 7012 6604 7064 6656
rect 7840 6672 7892 6724
rect 8668 6672 8720 6724
rect 10324 6672 10376 6724
rect 10508 6672 10560 6724
rect 7932 6604 7984 6656
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 12808 6672 12860 6724
rect 14096 6715 14148 6724
rect 13084 6604 13136 6656
rect 14096 6681 14105 6715
rect 14105 6681 14139 6715
rect 14139 6681 14148 6715
rect 14096 6672 14148 6681
rect 14188 6672 14240 6724
rect 18052 6740 18104 6792
rect 15752 6672 15804 6724
rect 15936 6672 15988 6724
rect 17868 6672 17920 6724
rect 20996 6808 21048 6860
rect 19984 6740 20036 6792
rect 23112 6876 23164 6928
rect 23296 6876 23348 6928
rect 25596 6876 25648 6928
rect 22100 6808 22152 6860
rect 22008 6740 22060 6792
rect 22284 6740 22336 6792
rect 22652 6740 22704 6792
rect 26240 6808 26292 6860
rect 26516 6808 26568 6860
rect 23572 6740 23624 6792
rect 24308 6740 24360 6792
rect 26884 6808 26936 6860
rect 27436 6740 27488 6792
rect 27804 6851 27856 6860
rect 27804 6817 27813 6851
rect 27813 6817 27847 6851
rect 27847 6817 27856 6851
rect 27804 6808 27856 6817
rect 28816 6808 28868 6860
rect 29184 6808 29236 6860
rect 30564 6808 30616 6860
rect 18420 6672 18472 6724
rect 20536 6672 20588 6724
rect 20720 6715 20772 6724
rect 20720 6681 20729 6715
rect 20729 6681 20763 6715
rect 20763 6681 20772 6715
rect 20720 6672 20772 6681
rect 22928 6672 22980 6724
rect 26884 6715 26936 6724
rect 13268 6604 13320 6656
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16212 6604 16264 6656
rect 16672 6604 16724 6656
rect 20352 6604 20404 6656
rect 22560 6647 22612 6656
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 26884 6681 26893 6715
rect 26893 6681 26927 6715
rect 26927 6681 26936 6715
rect 26884 6672 26936 6681
rect 26976 6604 27028 6656
rect 27804 6715 27856 6724
rect 27804 6681 27813 6715
rect 27813 6681 27847 6715
rect 27847 6681 27856 6715
rect 27804 6672 27856 6681
rect 28172 6740 28224 6792
rect 28540 6783 28592 6792
rect 28540 6749 28549 6783
rect 28549 6749 28583 6783
rect 28583 6749 28592 6783
rect 28540 6740 28592 6749
rect 30196 6740 30248 6792
rect 31944 6783 31996 6792
rect 31944 6749 31953 6783
rect 31953 6749 31987 6783
rect 31987 6749 31996 6783
rect 31944 6740 31996 6749
rect 34704 6783 34756 6792
rect 30748 6672 30800 6724
rect 31668 6672 31720 6724
rect 29276 6604 29328 6656
rect 31300 6604 31352 6656
rect 31852 6604 31904 6656
rect 32220 6715 32272 6724
rect 32220 6681 32254 6715
rect 32254 6681 32272 6715
rect 32220 6672 32272 6681
rect 33968 6672 34020 6724
rect 34704 6749 34713 6783
rect 34713 6749 34747 6783
rect 34747 6749 34756 6783
rect 34704 6740 34756 6749
rect 34796 6672 34848 6724
rect 36820 6740 36872 6792
rect 37188 6740 37240 6792
rect 33600 6604 33652 6656
rect 35900 6604 35952 6656
rect 37372 6604 37424 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 5816 6400 5868 6452
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 3700 6332 3752 6384
rect 3884 6332 3936 6384
rect 4068 6332 4120 6384
rect 3608 6264 3660 6316
rect 4712 6332 4764 6384
rect 4804 6332 4856 6384
rect 5356 6332 5408 6384
rect 6460 6332 6512 6384
rect 7840 6400 7892 6452
rect 7932 6400 7984 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 3884 6196 3936 6248
rect 4068 6196 4120 6248
rect 5724 6264 5776 6316
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7932 6264 7984 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 7656 6196 7708 6248
rect 7748 6196 7800 6248
rect 8944 6264 8996 6316
rect 8392 6196 8444 6248
rect 11244 6400 11296 6452
rect 11980 6400 12032 6452
rect 12808 6400 12860 6452
rect 13268 6400 13320 6452
rect 9588 6264 9640 6316
rect 9680 6264 9732 6316
rect 10692 6332 10744 6384
rect 10968 6332 11020 6384
rect 13360 6332 13412 6384
rect 14004 6332 14056 6384
rect 15108 6375 15160 6384
rect 15108 6341 15117 6375
rect 15117 6341 15151 6375
rect 15151 6341 15160 6375
rect 15108 6332 15160 6341
rect 15384 6400 15436 6452
rect 15844 6400 15896 6452
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 17224 6400 17276 6452
rect 17316 6400 17368 6452
rect 10232 6264 10284 6316
rect 12624 6264 12676 6316
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 14556 6264 14608 6316
rect 15016 6264 15068 6316
rect 15568 6332 15620 6384
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 17684 6332 17736 6384
rect 18604 6332 18656 6384
rect 19984 6443 20036 6452
rect 19984 6409 19993 6443
rect 19993 6409 20027 6443
rect 20027 6409 20036 6443
rect 19984 6400 20036 6409
rect 20444 6400 20496 6452
rect 20536 6400 20588 6452
rect 22468 6400 22520 6452
rect 22744 6400 22796 6452
rect 24032 6400 24084 6452
rect 24768 6400 24820 6452
rect 24860 6400 24912 6452
rect 26884 6400 26936 6452
rect 29736 6400 29788 6452
rect 31852 6400 31904 6452
rect 29276 6375 29328 6384
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 10968 6196 11020 6248
rect 12716 6196 12768 6248
rect 13084 6196 13136 6248
rect 19892 6264 19944 6316
rect 19984 6264 20036 6316
rect 20352 6264 20404 6316
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 21272 6264 21324 6316
rect 22100 6264 22152 6316
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 22652 6307 22704 6316
rect 22652 6273 22686 6307
rect 22686 6273 22704 6307
rect 22652 6264 22704 6273
rect 26056 6264 26108 6316
rect 26240 6264 26292 6316
rect 26700 6264 26752 6316
rect 29276 6341 29285 6375
rect 29285 6341 29319 6375
rect 29319 6341 29328 6375
rect 29276 6332 29328 6341
rect 29368 6332 29420 6384
rect 18052 6239 18104 6248
rect 3424 6060 3476 6112
rect 3700 6060 3752 6112
rect 8944 6128 8996 6180
rect 11152 6128 11204 6180
rect 5172 6060 5224 6112
rect 5448 6060 5500 6112
rect 6460 6060 6512 6112
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 6828 6060 6880 6112
rect 10324 6060 10376 6112
rect 10508 6060 10560 6112
rect 11796 6060 11848 6112
rect 12624 6128 12676 6180
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 23572 6196 23624 6248
rect 25320 6196 25372 6248
rect 15752 6128 15804 6180
rect 14832 6060 14884 6112
rect 15016 6060 15068 6112
rect 16672 6060 16724 6112
rect 17960 6060 18012 6112
rect 20444 6171 20496 6180
rect 20444 6137 20453 6171
rect 20453 6137 20487 6171
rect 20487 6137 20496 6171
rect 20444 6128 20496 6137
rect 24400 6128 24452 6180
rect 24032 6060 24084 6112
rect 24492 6103 24544 6112
rect 24492 6069 24501 6103
rect 24501 6069 24535 6103
rect 24535 6069 24544 6103
rect 24492 6060 24544 6069
rect 25136 6060 25188 6112
rect 25780 6103 25832 6112
rect 25780 6069 25789 6103
rect 25789 6069 25823 6103
rect 25823 6069 25832 6103
rect 25780 6060 25832 6069
rect 29644 6264 29696 6316
rect 30288 6264 30340 6316
rect 31116 6332 31168 6384
rect 32404 6375 32456 6384
rect 32404 6341 32413 6375
rect 32413 6341 32447 6375
rect 32447 6341 32456 6375
rect 32404 6332 32456 6341
rect 32588 6375 32640 6384
rect 32588 6341 32613 6375
rect 32613 6341 32640 6375
rect 32956 6400 33008 6452
rect 33416 6400 33468 6452
rect 34244 6400 34296 6452
rect 36176 6400 36228 6452
rect 32588 6332 32640 6341
rect 33232 6332 33284 6384
rect 34152 6332 34204 6384
rect 30472 6264 30524 6316
rect 31668 6264 31720 6316
rect 34796 6264 34848 6316
rect 35808 6332 35860 6384
rect 28080 6196 28132 6248
rect 30840 6196 30892 6248
rect 31208 6196 31260 6248
rect 32496 6128 32548 6180
rect 33416 6196 33468 6248
rect 34704 6196 34756 6248
rect 36820 6196 36872 6248
rect 34336 6128 34388 6180
rect 28172 6060 28224 6112
rect 28264 6060 28316 6112
rect 28724 6060 28776 6112
rect 29460 6103 29512 6112
rect 29460 6069 29469 6103
rect 29469 6069 29503 6103
rect 29503 6069 29512 6103
rect 29460 6060 29512 6069
rect 29736 6060 29788 6112
rect 30104 6060 30156 6112
rect 31024 6060 31076 6112
rect 33784 6060 33836 6112
rect 34428 6060 34480 6112
rect 36360 6060 36412 6112
rect 37464 6060 37516 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5540 5899 5592 5908
rect 3700 5788 3752 5840
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 10968 5856 11020 5908
rect 11336 5856 11388 5908
rect 11980 5856 12032 5908
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 14648 5856 14700 5908
rect 15016 5856 15068 5908
rect 15200 5856 15252 5908
rect 16120 5856 16172 5908
rect 20352 5856 20404 5908
rect 23388 5856 23440 5908
rect 23480 5899 23532 5908
rect 23480 5865 23489 5899
rect 23489 5865 23523 5899
rect 23523 5865 23532 5899
rect 23480 5856 23532 5865
rect 25320 5856 25372 5908
rect 26056 5856 26108 5908
rect 8668 5788 8720 5840
rect 8944 5788 8996 5840
rect 2504 5652 2556 5704
rect 3148 5720 3200 5772
rect 4068 5720 4120 5772
rect 5816 5720 5868 5772
rect 9128 5652 9180 5704
rect 5264 5584 5316 5636
rect 6092 5584 6144 5636
rect 7196 5584 7248 5636
rect 3884 5516 3936 5568
rect 5080 5516 5132 5568
rect 6920 5516 6972 5568
rect 8208 5627 8260 5636
rect 8208 5593 8217 5627
rect 8217 5593 8251 5627
rect 8251 5593 8260 5627
rect 8208 5584 8260 5593
rect 10232 5652 10284 5704
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 10048 5516 10100 5568
rect 12532 5720 12584 5772
rect 14188 5788 14240 5840
rect 14924 5788 14976 5840
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 15752 5788 15804 5840
rect 16948 5788 17000 5840
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 16120 5720 16172 5772
rect 14188 5584 14240 5636
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 14924 5584 14976 5636
rect 15384 5652 15436 5704
rect 16856 5720 16908 5772
rect 17224 5720 17276 5772
rect 16580 5652 16632 5704
rect 17592 5720 17644 5772
rect 17684 5652 17736 5704
rect 17960 5720 18012 5772
rect 18052 5720 18104 5772
rect 22744 5788 22796 5840
rect 27804 5856 27856 5908
rect 29460 5856 29512 5908
rect 31208 5856 31260 5908
rect 31760 5856 31812 5908
rect 33784 5899 33836 5908
rect 33784 5865 33793 5899
rect 33793 5865 33827 5899
rect 33827 5865 33836 5899
rect 33784 5856 33836 5865
rect 33876 5856 33928 5908
rect 34428 5856 34480 5908
rect 34612 5856 34664 5908
rect 36452 5856 36504 5908
rect 29368 5788 29420 5840
rect 30012 5788 30064 5840
rect 23572 5763 23624 5772
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 19340 5652 19392 5704
rect 15936 5584 15988 5636
rect 13636 5516 13688 5568
rect 17040 5516 17092 5568
rect 22008 5695 22060 5704
rect 22008 5661 22017 5695
rect 22017 5661 22051 5695
rect 22051 5661 22060 5695
rect 23572 5729 23581 5763
rect 23581 5729 23615 5763
rect 23615 5729 23624 5763
rect 23572 5720 23624 5729
rect 27436 5720 27488 5772
rect 30380 5788 30432 5840
rect 30288 5720 30340 5772
rect 32588 5720 32640 5772
rect 22008 5652 22060 5661
rect 22928 5652 22980 5704
rect 23388 5652 23440 5704
rect 24308 5652 24360 5704
rect 27528 5652 27580 5704
rect 27712 5652 27764 5704
rect 28816 5652 28868 5704
rect 29000 5695 29052 5704
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 29368 5652 29420 5704
rect 30748 5695 30800 5704
rect 24492 5584 24544 5636
rect 26884 5584 26936 5636
rect 26976 5584 27028 5636
rect 21732 5516 21784 5568
rect 22744 5516 22796 5568
rect 23296 5516 23348 5568
rect 23664 5516 23716 5568
rect 28724 5516 28776 5568
rect 29828 5584 29880 5636
rect 30748 5661 30757 5695
rect 30757 5661 30791 5695
rect 30791 5661 30800 5695
rect 30748 5652 30800 5661
rect 28908 5516 28960 5568
rect 31300 5584 31352 5636
rect 30380 5516 30432 5568
rect 32956 5627 33008 5636
rect 32956 5593 32981 5627
rect 32981 5593 33008 5627
rect 33232 5652 33284 5704
rect 36084 5652 36136 5704
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 33600 5627 33652 5636
rect 32956 5584 33008 5593
rect 33600 5593 33609 5627
rect 33609 5593 33643 5627
rect 33643 5593 33652 5627
rect 33600 5584 33652 5593
rect 36544 5584 36596 5636
rect 34796 5516 34848 5568
rect 35532 5516 35584 5568
rect 35992 5516 36044 5568
rect 37096 5559 37148 5568
rect 37096 5525 37105 5559
rect 37105 5525 37139 5559
rect 37139 5525 37148 5559
rect 37096 5516 37148 5525
rect 39396 5516 39448 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 4068 5244 4120 5296
rect 4620 5244 4672 5296
rect 4896 5312 4948 5364
rect 8116 5312 8168 5364
rect 9036 5312 9088 5364
rect 10140 5312 10192 5364
rect 10324 5312 10376 5364
rect 11980 5312 12032 5364
rect 13544 5312 13596 5364
rect 14096 5312 14148 5364
rect 3056 5176 3108 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 6460 5176 6512 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7380 5244 7432 5296
rect 8668 5244 8720 5296
rect 7472 5176 7524 5228
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9772 5244 9824 5296
rect 10876 5244 10928 5296
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 4068 4972 4120 5024
rect 10048 5108 10100 5160
rect 10968 5108 11020 5160
rect 4712 5040 4764 5092
rect 5724 5040 5776 5092
rect 8300 5040 8352 5092
rect 11152 5176 11204 5228
rect 11428 5176 11480 5228
rect 11612 5176 11664 5228
rect 12532 5219 12584 5228
rect 12532 5185 12548 5219
rect 12548 5185 12582 5219
rect 12582 5185 12584 5219
rect 12532 5176 12584 5185
rect 13084 5176 13136 5228
rect 15384 5244 15436 5296
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 19432 5312 19484 5364
rect 22560 5312 22612 5364
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16488 5176 16540 5228
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 13912 5108 13964 5160
rect 15292 5108 15344 5160
rect 15384 5108 15436 5160
rect 6092 4972 6144 5024
rect 6368 4972 6420 5024
rect 12532 5040 12584 5092
rect 15292 4972 15344 5024
rect 15476 4972 15528 5024
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 20812 5108 20864 5160
rect 22284 5176 22336 5228
rect 22744 5176 22796 5228
rect 23296 5176 23348 5228
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 24308 5219 24360 5228
rect 23664 5176 23716 5185
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 20444 5040 20496 5092
rect 24032 5108 24084 5160
rect 25320 5244 25372 5296
rect 27712 5244 27764 5296
rect 24952 5219 25004 5228
rect 24952 5185 24961 5219
rect 24961 5185 24995 5219
rect 24995 5185 25004 5219
rect 25596 5219 25648 5228
rect 24952 5176 25004 5185
rect 25596 5185 25605 5219
rect 25605 5185 25639 5219
rect 25639 5185 25648 5219
rect 25596 5176 25648 5185
rect 25688 5176 25740 5228
rect 28908 5312 28960 5364
rect 28540 5244 28592 5296
rect 29276 5244 29328 5296
rect 30472 5312 30524 5364
rect 29736 5176 29788 5228
rect 29920 5244 29972 5296
rect 31852 5312 31904 5364
rect 33048 5312 33100 5364
rect 33324 5355 33376 5364
rect 33324 5321 33333 5355
rect 33333 5321 33367 5355
rect 33367 5321 33376 5355
rect 33324 5312 33376 5321
rect 32128 5287 32180 5296
rect 32128 5253 32137 5287
rect 32137 5253 32171 5287
rect 32171 5253 32180 5287
rect 32128 5244 32180 5253
rect 32496 5244 32548 5296
rect 30840 5176 30892 5228
rect 17224 4972 17276 5024
rect 18696 4972 18748 5024
rect 19432 4972 19484 5024
rect 21364 4972 21416 5024
rect 22468 5040 22520 5092
rect 22652 5083 22704 5092
rect 22652 5049 22661 5083
rect 22661 5049 22695 5083
rect 22695 5049 22704 5083
rect 22652 5040 22704 5049
rect 22284 4972 22336 5024
rect 25320 5040 25372 5092
rect 23480 4972 23532 5024
rect 24768 5015 24820 5024
rect 24768 4981 24777 5015
rect 24777 4981 24811 5015
rect 24811 4981 24820 5015
rect 24768 4972 24820 4981
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 26056 5015 26108 5024
rect 26056 4981 26065 5015
rect 26065 4981 26099 5015
rect 26099 4981 26108 5015
rect 26056 4972 26108 4981
rect 26884 4972 26936 5024
rect 27068 4972 27120 5024
rect 27436 5108 27488 5160
rect 31944 5176 31996 5228
rect 36544 5312 36596 5364
rect 36268 5244 36320 5296
rect 38108 5312 38160 5364
rect 33968 5219 34020 5228
rect 33968 5185 33977 5219
rect 33977 5185 34011 5219
rect 34011 5185 34020 5219
rect 33968 5176 34020 5185
rect 36544 5176 36596 5228
rect 28632 5040 28684 5092
rect 28816 4972 28868 5024
rect 30196 5015 30248 5024
rect 30196 4981 30205 5015
rect 30205 4981 30239 5015
rect 30239 4981 30248 5015
rect 30196 4972 30248 4981
rect 34704 5108 34756 5160
rect 33232 5040 33284 5092
rect 34336 5040 34388 5092
rect 31668 4972 31720 5024
rect 31760 4972 31812 5024
rect 32588 4972 32640 5024
rect 34428 5015 34480 5024
rect 34428 4981 34437 5015
rect 34437 4981 34471 5015
rect 34471 4981 34480 5015
rect 34428 4972 34480 4981
rect 36452 4972 36504 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 3792 4768 3844 4820
rect 4804 4768 4856 4820
rect 5448 4768 5500 4820
rect 6920 4768 6972 4820
rect 7564 4768 7616 4820
rect 9312 4768 9364 4820
rect 5816 4700 5868 4752
rect 6368 4700 6420 4752
rect 8576 4700 8628 4752
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 6000 4632 6052 4684
rect 9772 4700 9824 4752
rect 4160 4564 4212 4616
rect 4344 4564 4396 4616
rect 4988 4564 5040 4616
rect 5448 4607 5500 4616
rect 5448 4573 5458 4607
rect 5458 4573 5492 4607
rect 5492 4573 5500 4607
rect 5448 4564 5500 4573
rect 5632 4564 5684 4616
rect 5908 4564 5960 4616
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 14556 4768 14608 4820
rect 15200 4768 15252 4820
rect 10508 4700 10560 4752
rect 6828 4564 6880 4616
rect 3792 4496 3844 4548
rect 4068 4539 4120 4548
rect 4068 4505 4077 4539
rect 4077 4505 4111 4539
rect 4111 4505 4120 4539
rect 4068 4496 4120 4505
rect 7932 4564 7984 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 10968 4700 11020 4752
rect 12164 4700 12216 4752
rect 12256 4700 12308 4752
rect 13084 4700 13136 4752
rect 9220 4564 9272 4573
rect 8024 4539 8076 4548
rect 2320 4428 2372 4480
rect 3240 4428 3292 4480
rect 3424 4428 3476 4480
rect 8024 4505 8033 4539
rect 8033 4505 8067 4539
rect 8067 4505 8076 4539
rect 8024 4496 8076 4505
rect 8668 4496 8720 4548
rect 9956 4496 10008 4548
rect 4252 4428 4304 4480
rect 11612 4564 11664 4616
rect 11980 4564 12032 4616
rect 14096 4632 14148 4684
rect 12348 4496 12400 4548
rect 11152 4428 11204 4480
rect 12256 4428 12308 4480
rect 12808 4428 12860 4480
rect 13452 4564 13504 4616
rect 16672 4700 16724 4752
rect 21272 4700 21324 4752
rect 14280 4632 14332 4684
rect 15568 4632 15620 4684
rect 25412 4768 25464 4820
rect 27068 4768 27120 4820
rect 28816 4811 28868 4820
rect 28816 4777 28825 4811
rect 28825 4777 28859 4811
rect 28859 4777 28868 4811
rect 28816 4768 28868 4777
rect 15108 4564 15160 4616
rect 15292 4564 15344 4616
rect 15016 4496 15068 4548
rect 20444 4564 20496 4616
rect 26056 4700 26108 4752
rect 30748 4768 30800 4820
rect 31760 4768 31812 4820
rect 32036 4768 32088 4820
rect 32588 4811 32640 4820
rect 32588 4777 32597 4811
rect 32597 4777 32631 4811
rect 32631 4777 32640 4811
rect 32588 4768 32640 4777
rect 22836 4607 22888 4616
rect 16672 4496 16724 4548
rect 16764 4539 16816 4548
rect 16764 4505 16773 4539
rect 16773 4505 16807 4539
rect 16807 4505 16816 4539
rect 17316 4539 17368 4548
rect 16764 4496 16816 4505
rect 17316 4505 17325 4539
rect 17325 4505 17359 4539
rect 17359 4505 17368 4539
rect 17316 4496 17368 4505
rect 18144 4539 18196 4548
rect 14280 4428 14332 4480
rect 14648 4428 14700 4480
rect 17684 4471 17736 4480
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 18144 4505 18153 4539
rect 18153 4505 18187 4539
rect 18187 4505 18196 4539
rect 18144 4496 18196 4505
rect 20352 4496 20404 4548
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 20812 4471 20864 4480
rect 20812 4437 20821 4471
rect 20821 4437 20855 4471
rect 20855 4437 20864 4471
rect 20812 4428 20864 4437
rect 20904 4428 20956 4480
rect 22284 4471 22336 4480
rect 22284 4437 22293 4471
rect 22293 4437 22327 4471
rect 22327 4437 22336 4471
rect 22284 4428 22336 4437
rect 22468 4428 22520 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24216 4428 24268 4480
rect 24676 4564 24728 4616
rect 26884 4607 26936 4616
rect 26884 4573 26893 4607
rect 26893 4573 26927 4607
rect 26927 4573 26936 4607
rect 26884 4564 26936 4573
rect 27160 4564 27212 4616
rect 24952 4496 25004 4548
rect 25320 4496 25372 4548
rect 26056 4496 26108 4548
rect 26516 4496 26568 4548
rect 27068 4496 27120 4548
rect 29828 4632 29880 4684
rect 32220 4700 32272 4752
rect 34612 4768 34664 4820
rect 35348 4768 35400 4820
rect 35808 4768 35860 4820
rect 36452 4768 36504 4820
rect 38016 4768 38068 4820
rect 29092 4564 29144 4616
rect 28908 4496 28960 4548
rect 28540 4428 28592 4480
rect 29828 4496 29880 4548
rect 31300 4496 31352 4548
rect 33968 4632 34020 4684
rect 36084 4632 36136 4684
rect 31668 4564 31720 4616
rect 29920 4471 29972 4480
rect 29920 4437 29929 4471
rect 29929 4437 29963 4471
rect 29963 4437 29972 4471
rect 29920 4428 29972 4437
rect 30288 4428 30340 4480
rect 31852 4428 31904 4480
rect 32496 4496 32548 4548
rect 33048 4496 33100 4548
rect 33416 4607 33468 4616
rect 33416 4573 33425 4607
rect 33425 4573 33459 4607
rect 33459 4573 33468 4607
rect 33416 4564 33468 4573
rect 33600 4564 33652 4616
rect 36544 4564 36596 4616
rect 37648 4564 37700 4616
rect 34796 4496 34848 4548
rect 34888 4539 34940 4548
rect 34888 4505 34913 4539
rect 34913 4505 34940 4539
rect 34888 4496 34940 4505
rect 32312 4428 32364 4480
rect 33232 4471 33284 4480
rect 33232 4437 33241 4471
rect 33241 4437 33275 4471
rect 33275 4437 33284 4471
rect 33232 4428 33284 4437
rect 33416 4428 33468 4480
rect 34244 4428 34296 4480
rect 36084 4496 36136 4548
rect 36176 4496 36228 4548
rect 37924 4428 37976 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2320 4224 2372 4276
rect 3424 4224 3476 4276
rect 4252 4224 4304 4276
rect 2872 4088 2924 4140
rect 3608 4088 3660 4140
rect 3884 4088 3936 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4712 4224 4764 4276
rect 7380 4224 7432 4276
rect 8024 4224 8076 4276
rect 8668 4224 8720 4276
rect 11704 4224 11756 4276
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 11980 4224 12032 4276
rect 13084 4224 13136 4276
rect 2320 4020 2372 4072
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5816 4131 5868 4140
rect 5540 4088 5592 4097
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7012 4156 7064 4208
rect 6736 4088 6788 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7380 4088 7432 4140
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 8576 4156 8628 4208
rect 9588 4156 9640 4208
rect 9680 4156 9732 4208
rect 10416 4156 10468 4208
rect 12808 4199 12860 4208
rect 5356 4020 5408 4072
rect 3424 3952 3476 4004
rect 3700 3952 3752 4004
rect 5448 3952 5500 4004
rect 7564 4020 7616 4072
rect 7840 4020 7892 4072
rect 8208 4020 8260 4072
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 12808 4165 12817 4199
rect 12817 4165 12851 4199
rect 12851 4165 12860 4199
rect 12808 4156 12860 4165
rect 13268 4156 13320 4208
rect 14280 4224 14332 4276
rect 15200 4224 15252 4276
rect 14648 4156 14700 4208
rect 13176 4131 13228 4140
rect 11704 4088 11756 4097
rect 9956 4020 10008 4072
rect 11612 4020 11664 4072
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 14188 4088 14240 4140
rect 14280 4088 14332 4140
rect 14924 4156 14976 4208
rect 5632 3952 5684 4004
rect 11980 3952 12032 4004
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6000 3884 6052 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7932 3927 7984 3936
rect 7932 3893 7941 3927
rect 7941 3893 7975 3927
rect 7975 3893 7984 3927
rect 7932 3884 7984 3893
rect 8576 3884 8628 3936
rect 8944 3884 8996 3936
rect 11152 3884 11204 3936
rect 11336 3884 11388 3936
rect 11888 3884 11940 3936
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 14556 3952 14608 4004
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 16304 4224 16356 4276
rect 18052 4224 18104 4276
rect 20444 4267 20496 4276
rect 19616 4156 19668 4208
rect 20444 4233 20453 4267
rect 20453 4233 20487 4267
rect 20487 4233 20496 4267
rect 20444 4224 20496 4233
rect 22560 4224 22612 4276
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 17224 4088 17276 4140
rect 18880 4131 18932 4140
rect 18880 4097 18914 4131
rect 18914 4097 18932 4131
rect 18880 4088 18932 4097
rect 19156 4088 19208 4140
rect 19248 4088 19300 4140
rect 20168 4088 20220 4140
rect 21272 4156 21324 4208
rect 24032 4156 24084 4208
rect 24492 4156 24544 4208
rect 27436 4224 27488 4276
rect 29460 4224 29512 4276
rect 29920 4224 29972 4276
rect 30196 4224 30248 4276
rect 33232 4224 33284 4276
rect 34612 4224 34664 4276
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20996 4131 21048 4140
rect 20720 4088 20772 4097
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 22376 4088 22428 4140
rect 23480 4088 23532 4140
rect 24400 4131 24452 4140
rect 24400 4097 24409 4131
rect 24409 4097 24443 4131
rect 24443 4097 24452 4131
rect 24400 4088 24452 4097
rect 24676 4088 24728 4140
rect 24768 4088 24820 4140
rect 25688 4088 25740 4140
rect 25872 4088 25924 4140
rect 26424 4131 26476 4140
rect 26424 4097 26433 4131
rect 26433 4097 26467 4131
rect 26467 4097 26476 4131
rect 26424 4088 26476 4097
rect 26884 4088 26936 4140
rect 27344 4088 27396 4140
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 29092 4156 29144 4208
rect 29828 4156 29880 4208
rect 28816 4088 28868 4140
rect 30012 4131 30064 4140
rect 30012 4097 30021 4131
rect 30021 4097 30055 4131
rect 30055 4097 30064 4131
rect 30012 4088 30064 4097
rect 30288 4131 30340 4140
rect 30288 4097 30322 4131
rect 30322 4097 30340 4131
rect 30288 4088 30340 4097
rect 32312 4131 32364 4140
rect 32312 4097 32321 4131
rect 32321 4097 32355 4131
rect 32355 4097 32364 4131
rect 32496 4131 32548 4140
rect 32312 4088 32364 4097
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 35440 4156 35492 4208
rect 33324 4088 33376 4140
rect 34520 4088 34572 4140
rect 36728 4088 36780 4140
rect 37280 4131 37332 4140
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 16212 4020 16264 4072
rect 18236 4020 18288 4072
rect 18604 4063 18656 4072
rect 18604 4029 18613 4063
rect 18613 4029 18647 4063
rect 18647 4029 18656 4063
rect 18604 4020 18656 4029
rect 19708 4020 19760 4072
rect 26516 4020 26568 4072
rect 32128 4020 32180 4072
rect 15660 3952 15712 4004
rect 23296 3952 23348 4004
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 17040 3884 17092 3936
rect 19800 3884 19852 3936
rect 20168 3884 20220 3936
rect 23480 3884 23532 3936
rect 24952 3884 25004 3936
rect 26884 3884 26936 3936
rect 33416 3952 33468 4004
rect 31300 3884 31352 3936
rect 31484 3884 31536 3936
rect 37188 4020 37240 4072
rect 38660 3952 38712 4004
rect 34704 3884 34756 3936
rect 34796 3884 34848 3936
rect 35440 3884 35492 3936
rect 37188 3884 37240 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3332 3680 3384 3732
rect 6736 3680 6788 3732
rect 7288 3680 7340 3732
rect 12256 3680 12308 3732
rect 13268 3680 13320 3732
rect 15384 3680 15436 3732
rect 16948 3680 17000 3732
rect 5540 3612 5592 3664
rect 8116 3612 8168 3664
rect 8944 3612 8996 3664
rect 3700 3544 3752 3596
rect 7380 3544 7432 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 3240 3519 3292 3528
rect 1952 3476 2004 3485
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 4620 3476 4672 3528
rect 6736 3476 6788 3528
rect 8576 3544 8628 3596
rect 8852 3544 8904 3596
rect 5724 3408 5776 3460
rect 3884 3340 3936 3392
rect 7288 3340 7340 3392
rect 7380 3340 7432 3392
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 8116 3519 8168 3528
rect 7840 3476 7892 3485
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 12072 3612 12124 3664
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15108 3544 15160 3596
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 17316 3680 17368 3732
rect 18328 3680 18380 3732
rect 18788 3680 18840 3732
rect 18972 3680 19024 3732
rect 19340 3680 19392 3732
rect 19708 3680 19760 3732
rect 11244 3519 11296 3528
rect 11244 3485 11278 3519
rect 11278 3485 11296 3519
rect 9036 3408 9088 3460
rect 9312 3408 9364 3460
rect 11244 3476 11296 3485
rect 12440 3476 12492 3528
rect 12532 3476 12584 3528
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 13268 3476 13320 3528
rect 14096 3476 14148 3528
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14648 3519 14700 3528
rect 14372 3476 14424 3485
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 15200 3476 15252 3528
rect 18236 3544 18288 3596
rect 18604 3612 18656 3664
rect 9588 3340 9640 3392
rect 9680 3340 9732 3392
rect 10324 3340 10376 3392
rect 11520 3408 11572 3460
rect 13176 3451 13228 3460
rect 13176 3417 13185 3451
rect 13185 3417 13219 3451
rect 13219 3417 13228 3451
rect 13176 3408 13228 3417
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 14832 3408 14884 3460
rect 15384 3408 15436 3460
rect 17408 3340 17460 3392
rect 18236 3408 18288 3460
rect 19064 3408 19116 3460
rect 20352 3544 20404 3596
rect 22376 3680 22428 3732
rect 26240 3680 26292 3732
rect 29000 3680 29052 3732
rect 32496 3680 32548 3732
rect 33968 3723 34020 3732
rect 33968 3689 33977 3723
rect 33977 3689 34011 3723
rect 34011 3689 34020 3723
rect 33968 3680 34020 3689
rect 34152 3723 34204 3732
rect 34152 3689 34161 3723
rect 34161 3689 34195 3723
rect 34195 3689 34204 3723
rect 34152 3680 34204 3689
rect 23112 3612 23164 3664
rect 23756 3612 23808 3664
rect 19892 3476 19944 3528
rect 19524 3408 19576 3460
rect 20168 3340 20220 3392
rect 20536 3476 20588 3528
rect 23388 3544 23440 3596
rect 20720 3476 20772 3528
rect 20996 3476 21048 3528
rect 23020 3519 23072 3528
rect 20812 3408 20864 3460
rect 21180 3451 21232 3460
rect 21180 3417 21214 3451
rect 21214 3417 21232 3451
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 21180 3408 21232 3417
rect 23480 3408 23532 3460
rect 21456 3340 21508 3392
rect 23296 3340 23348 3392
rect 26516 3655 26568 3664
rect 26516 3621 26525 3655
rect 26525 3621 26559 3655
rect 26559 3621 26568 3655
rect 26516 3612 26568 3621
rect 28908 3612 28960 3664
rect 34336 3612 34388 3664
rect 35440 3680 35492 3732
rect 36084 3723 36136 3732
rect 36084 3689 36093 3723
rect 36093 3689 36127 3723
rect 36127 3689 36136 3723
rect 36084 3680 36136 3689
rect 36912 3723 36964 3732
rect 36912 3689 36921 3723
rect 36921 3689 36955 3723
rect 36955 3689 36964 3723
rect 36912 3680 36964 3689
rect 36452 3612 36504 3664
rect 25872 3544 25924 3596
rect 26056 3544 26108 3596
rect 27252 3544 27304 3596
rect 27712 3544 27764 3596
rect 28724 3544 28776 3596
rect 29828 3587 29880 3596
rect 24216 3476 24268 3528
rect 26608 3476 26660 3528
rect 26884 3476 26936 3528
rect 27620 3408 27672 3460
rect 27804 3476 27856 3528
rect 28264 3476 28316 3528
rect 28632 3519 28684 3528
rect 28632 3485 28641 3519
rect 28641 3485 28675 3519
rect 28675 3485 28684 3519
rect 28632 3476 28684 3485
rect 29828 3553 29837 3587
rect 29837 3553 29871 3587
rect 29871 3553 29880 3587
rect 29828 3544 29880 3553
rect 30012 3544 30064 3596
rect 29736 3476 29788 3528
rect 30196 3476 30248 3528
rect 32864 3544 32916 3596
rect 34704 3587 34756 3596
rect 32128 3476 32180 3528
rect 32312 3476 32364 3528
rect 33324 3519 33376 3528
rect 33324 3485 33333 3519
rect 33333 3485 33367 3519
rect 33367 3485 33376 3519
rect 33324 3476 33376 3485
rect 34704 3553 34713 3587
rect 34713 3553 34747 3587
rect 34747 3553 34756 3587
rect 34704 3544 34756 3553
rect 31116 3408 31168 3460
rect 31484 3408 31536 3460
rect 33508 3408 33560 3460
rect 34612 3476 34664 3528
rect 37372 3519 37424 3528
rect 37372 3485 37381 3519
rect 37381 3485 37415 3519
rect 37415 3485 37424 3519
rect 37372 3476 37424 3485
rect 35624 3408 35676 3460
rect 36084 3408 36136 3460
rect 24032 3340 24084 3392
rect 24124 3340 24176 3392
rect 27252 3340 27304 3392
rect 27896 3340 27948 3392
rect 28448 3383 28500 3392
rect 28448 3349 28457 3383
rect 28457 3349 28491 3383
rect 28491 3349 28500 3383
rect 28448 3340 28500 3349
rect 29092 3340 29144 3392
rect 32864 3383 32916 3392
rect 32864 3349 32873 3383
rect 32873 3349 32907 3383
rect 32907 3349 32916 3383
rect 32864 3340 32916 3349
rect 36728 3383 36780 3392
rect 36728 3349 36753 3383
rect 36753 3349 36780 3383
rect 36728 3340 36780 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 3148 3136 3200 3188
rect 3240 3136 3292 3188
rect 4068 3136 4120 3188
rect 3608 3111 3660 3120
rect 3608 3077 3617 3111
rect 3617 3077 3651 3111
rect 3651 3077 3660 3111
rect 3608 3068 3660 3077
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 2780 3000 2832 3052
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4988 3136 5040 3188
rect 6828 3136 6880 3188
rect 5172 3000 5224 3052
rect 6368 3068 6420 3120
rect 8024 3136 8076 3188
rect 8484 3136 8536 3188
rect 8576 3136 8628 3188
rect 7196 3068 7248 3120
rect 5540 3000 5592 3052
rect 6092 3000 6144 3052
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 6552 2932 6604 2984
rect 7564 3000 7616 3052
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 9128 3043 9180 3052
rect 8852 3000 8904 3009
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 9496 2932 9548 2984
rect 11612 3000 11664 3052
rect 11980 3000 12032 3052
rect 11520 2975 11572 2984
rect 3608 2864 3660 2916
rect 5632 2796 5684 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 8116 2796 8168 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 9220 2796 9272 2848
rect 9404 2796 9456 2848
rect 10784 2864 10836 2916
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 12440 3000 12492 3052
rect 12256 2932 12308 2984
rect 14924 3136 14976 3188
rect 16856 3136 16908 3188
rect 19432 3136 19484 3188
rect 15844 3068 15896 3120
rect 15384 3000 15436 3052
rect 16028 3000 16080 3052
rect 18052 3068 18104 3120
rect 19248 3000 19300 3052
rect 19800 3000 19852 3052
rect 20812 3136 20864 3188
rect 20352 3068 20404 3120
rect 24308 3136 24360 3188
rect 25596 3136 25648 3188
rect 26148 3179 26200 3188
rect 26148 3145 26157 3179
rect 26157 3145 26191 3179
rect 26191 3145 26200 3179
rect 26148 3136 26200 3145
rect 29092 3179 29144 3188
rect 29092 3145 29101 3179
rect 29101 3145 29135 3179
rect 29135 3145 29144 3179
rect 29092 3136 29144 3145
rect 24032 3068 24084 3120
rect 20444 3000 20496 3052
rect 20536 3000 20588 3052
rect 21456 3000 21508 3052
rect 12164 2864 12216 2916
rect 14372 2864 14424 2916
rect 11796 2796 11848 2848
rect 12440 2796 12492 2848
rect 21088 2932 21140 2984
rect 23388 3000 23440 3052
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 24768 3000 24820 3052
rect 23480 2975 23532 2984
rect 23480 2941 23489 2975
rect 23489 2941 23523 2975
rect 23523 2941 23532 2975
rect 23480 2932 23532 2941
rect 24216 2932 24268 2984
rect 25228 3000 25280 3052
rect 25964 3043 26016 3052
rect 25964 3009 25973 3043
rect 25973 3009 26007 3043
rect 26007 3009 26016 3043
rect 25964 3000 26016 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 28172 3068 28224 3120
rect 30012 3136 30064 3188
rect 33508 3179 33560 3188
rect 33508 3145 33517 3179
rect 33517 3145 33551 3179
rect 33551 3145 33560 3179
rect 33508 3136 33560 3145
rect 34612 3136 34664 3188
rect 27804 3000 27856 3052
rect 28448 3000 28500 3052
rect 28908 3000 28960 3052
rect 32220 3068 32272 3120
rect 32864 3068 32916 3120
rect 34796 3111 34848 3120
rect 34796 3077 34805 3111
rect 34805 3077 34839 3111
rect 34839 3077 34848 3111
rect 34796 3068 34848 3077
rect 31944 3000 31996 3052
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 25872 2932 25924 2984
rect 28724 2932 28776 2984
rect 31392 2932 31444 2984
rect 33600 3000 33652 3052
rect 33692 3000 33744 3052
rect 35900 3068 35952 3120
rect 36636 3136 36688 3188
rect 36820 3068 36872 3120
rect 36728 3000 36780 3052
rect 37464 3000 37516 3052
rect 18328 2864 18380 2916
rect 16120 2796 16172 2848
rect 18236 2796 18288 2848
rect 18880 2839 18932 2848
rect 18880 2805 18889 2839
rect 18889 2805 18923 2839
rect 18923 2805 18932 2839
rect 18880 2796 18932 2805
rect 19340 2839 19392 2848
rect 19340 2805 19349 2839
rect 19349 2805 19383 2839
rect 19383 2805 19392 2839
rect 19340 2796 19392 2805
rect 19616 2796 19668 2848
rect 22744 2864 22796 2916
rect 20996 2796 21048 2848
rect 21640 2796 21692 2848
rect 22284 2796 22336 2848
rect 24308 2839 24360 2848
rect 24308 2805 24317 2839
rect 24317 2805 24351 2839
rect 24351 2805 24360 2839
rect 24308 2796 24360 2805
rect 25320 2864 25372 2916
rect 27712 2864 27764 2916
rect 29092 2864 29144 2916
rect 27620 2796 27672 2848
rect 29000 2796 29052 2848
rect 29736 2839 29788 2848
rect 29736 2805 29745 2839
rect 29745 2805 29779 2839
rect 29779 2805 29788 2839
rect 29736 2796 29788 2805
rect 35716 2864 35768 2916
rect 32772 2796 32824 2848
rect 34336 2796 34388 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2964 2592 3016 2644
rect 5540 2592 5592 2644
rect 5724 2592 5776 2644
rect 6828 2592 6880 2644
rect 9036 2592 9088 2644
rect 10416 2592 10468 2644
rect 12440 2592 12492 2644
rect 2688 2524 2740 2576
rect 3884 2456 3936 2508
rect 12256 2524 12308 2576
rect 13820 2592 13872 2644
rect 15200 2592 15252 2644
rect 15936 2592 15988 2644
rect 17684 2592 17736 2644
rect 18144 2592 18196 2644
rect 18604 2592 18656 2644
rect 18788 2592 18840 2644
rect 20076 2592 20128 2644
rect 20628 2592 20680 2644
rect 6828 2456 6880 2508
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 9404 2456 9456 2508
rect 8576 2388 8628 2440
rect 9956 2388 10008 2440
rect 10508 2431 10560 2440
rect 572 2320 624 2372
rect 7288 2320 7340 2372
rect 8484 2320 8536 2372
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 13820 2456 13872 2508
rect 15016 2456 15068 2508
rect 17224 2524 17276 2576
rect 17500 2524 17552 2576
rect 19340 2524 19392 2576
rect 15568 2456 15620 2508
rect 12992 2388 13044 2440
rect 16672 2456 16724 2508
rect 18788 2456 18840 2508
rect 24584 2524 24636 2576
rect 10876 2320 10928 2372
rect 14096 2320 14148 2372
rect 3148 2252 3200 2304
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 13268 2295 13320 2304
rect 13268 2261 13277 2295
rect 13277 2261 13311 2295
rect 13311 2261 13320 2295
rect 13268 2252 13320 2261
rect 16212 2388 16264 2440
rect 18052 2388 18104 2440
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18604 2431 18656 2440
rect 18328 2388 18380 2397
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 18880 2388 18932 2440
rect 19524 2388 19576 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 23296 2456 23348 2508
rect 24768 2499 24820 2508
rect 24768 2465 24777 2499
rect 24777 2465 24811 2499
rect 24811 2465 24820 2499
rect 24768 2456 24820 2465
rect 27068 2456 27120 2508
rect 29000 2592 29052 2644
rect 32036 2592 32088 2644
rect 30564 2524 30616 2576
rect 33508 2524 33560 2576
rect 34980 2524 35032 2576
rect 22008 2388 22060 2440
rect 22192 2388 22244 2440
rect 24860 2388 24912 2440
rect 15936 2252 15988 2304
rect 16488 2252 16540 2304
rect 24308 2320 24360 2372
rect 25504 2388 25556 2440
rect 26424 2388 26476 2440
rect 30840 2456 30892 2508
rect 28356 2388 28408 2440
rect 30380 2388 30432 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 34428 2456 34480 2508
rect 26240 2320 26292 2372
rect 26884 2320 26936 2372
rect 33140 2388 33192 2440
rect 35992 2456 36044 2508
rect 37096 2456 37148 2508
rect 36360 2388 36412 2440
rect 20628 2252 20680 2304
rect 23848 2252 23900 2304
rect 26056 2252 26108 2304
rect 35532 2320 35584 2372
rect 39764 2320 39816 2372
rect 29828 2252 29880 2304
rect 31300 2252 31352 2304
rect 34244 2252 34296 2304
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3332 2048 3384 2100
rect 4620 2048 4672 2100
rect 5172 2048 5224 2100
rect 13268 2048 13320 2100
rect 16396 2048 16448 2100
rect 22192 2048 22244 2100
rect 2504 1980 2556 2032
rect 9404 1980 9456 2032
rect 12256 1980 12308 2032
rect 3792 1912 3844 1964
rect 3056 1844 3108 1896
rect 10508 1844 10560 1896
rect 2412 1776 2464 1828
rect 7196 1776 7248 1828
rect 18604 1980 18656 2032
rect 30932 2048 30984 2100
rect 19800 1912 19852 1964
rect 21272 1912 21324 1964
rect 21456 1912 21508 1964
rect 38016 1980 38068 2032
rect 20444 1844 20496 1896
rect 21364 1776 21416 1828
rect 18328 1708 18380 1760
rect 22100 1708 22152 1760
rect 3976 1504 4028 1556
rect 5356 1504 5408 1556
rect 1860 1368 1912 1420
rect 7932 1368 7984 1420
rect 17960 1368 18012 1420
rect 20628 1368 20680 1420
rect 28356 1368 28408 1420
rect 29828 1368 29880 1420
rect 2780 1232 2832 1284
rect 4252 1232 4304 1284
rect 2596 1096 2648 1148
rect 9036 1096 9088 1148
<< metal2 >>
rect 4986 49314 5042 50000
rect 14922 49314 14978 50000
rect 24950 49314 25006 50000
rect 34978 49314 35034 50000
rect 4986 49286 5120 49314
rect 4986 49200 5042 49286
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 5092 47054 5120 49286
rect 14922 49286 15148 49314
rect 14922 49200 14978 49286
rect 15120 48090 15148 49286
rect 24950 49286 25268 49314
rect 24950 49200 25006 49286
rect 15120 48062 15240 48090
rect 15212 47258 15240 48062
rect 25240 47258 25268 49286
rect 34978 49286 35388 49314
rect 34978 49200 35034 49286
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35360 47258 35388 49286
rect 15200 47252 15252 47258
rect 15200 47194 15252 47200
rect 25228 47252 25280 47258
rect 25228 47194 25280 47200
rect 35348 47252 35400 47258
rect 35348 47194 35400 47200
rect 5080 47048 5132 47054
rect 5080 46990 5132 46996
rect 19248 47048 19300 47054
rect 19248 46990 19300 46996
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 35348 47048 35400 47054
rect 35348 46990 35400 46996
rect 5264 46912 5316 46918
rect 5264 46854 5316 46860
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 5276 25362 5304 46854
rect 19260 46714 19288 46990
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19248 46708 19300 46714
rect 19248 46650 19300 46656
rect 20536 46572 20588 46578
rect 20536 46514 20588 46520
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19260 30326 19288 30534
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 15764 29714 15792 30194
rect 18432 29850 18460 30194
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 15752 29708 15804 29714
rect 15752 29650 15804 29656
rect 15764 28626 15792 29650
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16684 29306 16712 29514
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15384 28076 15436 28082
rect 15436 28036 15516 28064
rect 15384 28018 15436 28024
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 15304 27402 15332 27950
rect 15488 27538 15516 28036
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12452 26382 12480 27270
rect 13372 27130 13400 27338
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14200 26586 14228 26930
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 11808 23730 11836 25774
rect 12268 25498 12296 25842
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12360 23798 12388 24006
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 11808 22642 11836 23666
rect 12452 23186 12480 26318
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24886 12848 25094
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 13096 24818 13124 26250
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 13188 25294 13216 26182
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13176 25152 13228 25158
rect 13280 25106 13308 25638
rect 13228 25100 13308 25106
rect 13176 25094 13308 25100
rect 13188 25078 13308 25094
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13096 24206 13124 24754
rect 13188 24732 13216 25078
rect 13268 24744 13320 24750
rect 13188 24704 13268 24732
rect 13268 24686 13320 24692
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12544 23322 12572 24142
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 12452 22166 12480 23122
rect 12912 23118 12940 24006
rect 13096 23118 13124 24142
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13188 23866 13216 24074
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13096 22710 13124 22918
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 12820 21554 12848 22646
rect 13188 22522 13216 22918
rect 13096 22494 13216 22522
rect 13096 22030 13124 22494
rect 13280 22094 13308 24686
rect 13648 24682 13676 26318
rect 14936 26314 14964 27270
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14476 26042 14504 26250
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14752 25294 14780 25910
rect 14936 25906 14964 26250
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 14648 24744 14700 24750
rect 14752 24732 14780 25230
rect 14700 24704 14780 24732
rect 14648 24686 14700 24692
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24206 13400 24550
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13372 23118 13400 24142
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 13464 23594 13492 24074
rect 14660 23594 14688 24686
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13188 22066 13308 22094
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 12820 20602 12848 21490
rect 13096 21146 13124 21490
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 17270 10640 17546
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 10704 16454 10732 18226
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17202 11008 17478
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11072 17066 11100 18634
rect 11440 17746 11468 18702
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11256 16590 11284 17002
rect 11532 16658 11560 18158
rect 11808 17882 11836 18566
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11624 17270 11652 17546
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11716 16998 11744 17478
rect 11900 17338 11928 19314
rect 12636 19174 12664 20402
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12084 17678 12112 19110
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 12544 16998 12572 18022
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9508 15026 9536 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15162 9720 15302
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 10244 15094 10272 15846
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 9508 14482 9536 14962
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 9508 13326 9536 13806
rect 9784 13326 9812 14010
rect 10520 14006 10548 15506
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11830 8984 12038
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 6552 11688 6604 11694
rect 8484 11688 8536 11694
rect 6552 11630 6604 11636
rect 8404 11636 8484 11642
rect 8404 11630 8536 11636
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1596 8634 1624 10474
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4908 9654 4936 11086
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 5000 9586 5028 9862
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3988 9081 4016 9114
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8634 3464 8774
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3252 8537 3280 8570
rect 3238 8528 3294 8537
rect 3238 8463 3294 8472
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 8401 3648 8434
rect 3606 8392 3662 8401
rect 3606 8327 3662 8336
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 202 3360 258 3369
rect 202 3295 258 3304
rect 216 800 244 3295
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 584 800 612 2314
rect 952 800 980 7346
rect 1320 800 1348 7822
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 2318 7712 2374 7721
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1674 6488 1730 6497
rect 1674 6423 1676 6432
rect 1728 6423 1730 6432
rect 1676 6394 1728 6400
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 3097 1716 4966
rect 1780 3534 1808 7142
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1872 5137 1900 5170
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1964 3534 1992 7686
rect 2318 7647 2374 7656
rect 2332 7002 2360 7647
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4282 2360 4422
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 2332 3194 2360 4014
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1674 3088 1730 3097
rect 1674 3023 1730 3032
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 1426 1900 2994
rect 2424 1834 2452 6734
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5545 2544 5646
rect 2502 5536 2558 5545
rect 2502 5471 2558 5480
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 2038 2544 5170
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2504 2032 2556 2038
rect 2504 1974 2556 1980
rect 2412 1828 2464 1834
rect 2412 1770 2464 1776
rect 1860 1420 1912 1426
rect 1860 1362 1912 1368
rect 2608 1154 2636 4558
rect 2792 4162 2820 6734
rect 2884 4298 2912 7822
rect 2976 7002 3004 8230
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3238 7440 3294 7449
rect 3238 7375 3240 7384
rect 3292 7375 3294 7384
rect 3240 7346 3292 7352
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 7002 3096 7142
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2976 4434 3004 6394
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3160 5409 3188 5714
rect 3146 5400 3202 5409
rect 3146 5335 3202 5344
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 4826 3096 5170
rect 3056 4820 3108 4826
rect 3252 4808 3280 6734
rect 3056 4762 3108 4768
rect 3160 4780 3280 4808
rect 2976 4406 3096 4434
rect 2884 4270 3004 4298
rect 2700 4134 2820 4162
rect 2870 4176 2926 4185
rect 2700 2582 2728 4134
rect 2870 4111 2872 4120
rect 2924 4111 2926 4120
rect 2872 4082 2924 4088
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2792 1290 2820 2994
rect 2976 2650 3004 4270
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 1902 3096 4406
rect 3160 3618 3188 4780
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3252 4486 3280 4655
rect 3240 4480 3292 4486
rect 3344 4457 3372 7686
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5273 3464 6054
rect 3422 5264 3478 5273
rect 3422 5199 3478 5208
rect 3424 4480 3476 4486
rect 3240 4422 3292 4428
rect 3330 4448 3386 4457
rect 3424 4422 3476 4428
rect 3330 4383 3386 4392
rect 3436 4282 3464 4422
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3330 4176 3386 4185
rect 3330 4111 3386 4120
rect 3344 3738 3372 4111
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3641 3464 3946
rect 3422 3632 3478 3641
rect 3160 3590 3372 3618
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3146 3224 3202 3233
rect 3252 3194 3280 3470
rect 3146 3159 3148 3168
rect 3200 3159 3202 3168
rect 3240 3188 3292 3194
rect 3148 3130 3200 3136
rect 3240 3130 3292 3136
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3160 2961 3188 2994
rect 3146 2952 3202 2961
rect 3146 2887 3202 2896
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 2780 1284 2832 1290
rect 2780 1226 2832 1232
rect 2596 1148 2648 1154
rect 2596 1090 2648 1096
rect 3160 800 3188 2246
rect 3344 2106 3372 3590
rect 3422 3567 3478 3576
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3528 800 3556 7822
rect 3698 7576 3754 7585
rect 3698 7511 3700 7520
rect 3752 7511 3754 7520
rect 3700 7482 3752 7488
rect 3700 6384 3752 6390
rect 3698 6352 3700 6361
rect 3752 6352 3754 6361
rect 3608 6316 3660 6322
rect 3698 6287 3754 6296
rect 3608 6258 3660 6264
rect 3620 4264 3648 6258
rect 3698 6216 3754 6225
rect 3698 6151 3754 6160
rect 3712 6118 3740 6151
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3712 5681 3740 5782
rect 3698 5672 3754 5681
rect 3698 5607 3754 5616
rect 3804 4826 3832 8298
rect 3896 6866 3924 8910
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 4172 8809 4200 8842
rect 4158 8800 4214 8809
rect 4158 8735 4214 8744
rect 4066 8664 4122 8673
rect 4066 8599 4068 8608
rect 4120 8599 4122 8608
rect 4068 8570 4120 8576
rect 4724 8362 4752 8842
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4908 8090 4936 8434
rect 5078 8120 5134 8129
rect 4896 8084 4948 8090
rect 5078 8055 5134 8064
rect 4896 8026 4948 8032
rect 5092 7954 5120 8055
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4528 7880 4580 7886
rect 4526 7848 4528 7857
rect 4580 7848 4582 7857
rect 4526 7783 4582 7792
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 3976 7336 4028 7342
rect 4448 7313 4476 7346
rect 3976 7278 4028 7284
rect 4434 7304 4490 7313
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3896 6390 3924 6802
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5574 3924 6190
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3790 4584 3846 4593
rect 3790 4519 3792 4528
rect 3844 4519 3846 4528
rect 3792 4490 3844 4496
rect 3620 4236 3832 4264
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 4049 3648 4082
rect 3606 4040 3662 4049
rect 3606 3975 3662 3984
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3712 3602 3740 3946
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3804 3505 3832 4236
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3896 3398 3924 4082
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3620 2922 3648 3062
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3804 1970 3832 2382
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3896 800 3924 2450
rect 3988 1562 4016 7278
rect 4434 7239 4490 7248
rect 4896 7200 4948 7206
rect 4894 7168 4896 7177
rect 4948 7168 4950 7177
rect 4214 7100 4522 7120
rect 4894 7103 4950 7112
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6390 4108 6598
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4068 6248 4120 6254
rect 4540 6236 4568 6870
rect 4724 6390 4752 6870
rect 4804 6792 4856 6798
rect 4856 6752 5028 6780
rect 4804 6734 4856 6740
rect 5000 6662 5028 6752
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4816 6236 4844 6326
rect 4540 6208 4844 6236
rect 4068 6190 4120 6196
rect 4080 5778 4108 6190
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5302 4108 5714
rect 4908 5370 4936 6598
rect 5092 6089 5120 7686
rect 5184 7274 5212 8842
rect 5276 8566 5304 10134
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5368 8294 5396 9522
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8430 5580 9318
rect 5644 8894 5856 8922
rect 5644 8498 5672 8894
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 7936 5488 8298
rect 5460 7908 5672 7936
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5368 7721 5396 7754
rect 5354 7712 5410 7721
rect 5354 7647 5410 7656
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5368 6905 5396 7346
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5172 6112 5224 6118
rect 5078 6080 5134 6089
rect 5172 6054 5224 6060
rect 5078 6015 5134 6024
rect 4986 5808 5042 5817
rect 4986 5743 5042 5752
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4894 5264 4950 5273
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4554 4108 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 3194 4108 4490
rect 4172 4146 4200 4558
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4282 4292 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4356 4146 4384 4558
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3534 4660 5238
rect 4804 5228 4856 5234
rect 4894 5199 4950 5208
rect 4804 5170 4856 5176
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4282 4752 5034
rect 4816 4826 4844 5170
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4908 3913 4936 5199
rect 5000 4622 5028 5743
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4894 3904 4950 3913
rect 4894 3839 4950 3848
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5000 3194 5028 4558
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5092 2774 5120 5510
rect 5184 3058 5212 6054
rect 5368 5658 5396 6326
rect 5460 6118 5488 6802
rect 5552 6730 5580 7210
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5644 6610 5672 7908
rect 5736 7886 5764 8774
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5552 6582 5672 6610
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5552 5914 5580 6582
rect 5828 6458 5856 8894
rect 5920 6730 5948 9590
rect 6012 8129 6040 9862
rect 6288 9586 6316 11494
rect 6564 11150 6592 11630
rect 8404 11614 8524 11630
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6656 10810 6684 11018
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6564 9586 6592 10202
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9586 6684 9998
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8498 6132 8774
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5998 8120 6054 8129
rect 5998 8055 6000 8064
rect 6052 8055 6054 8064
rect 6000 8026 6052 8032
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5264 5636 5316 5642
rect 5368 5630 5488 5658
rect 5264 5578 5316 5584
rect 5276 4146 5304 5578
rect 5460 4826 5488 5630
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4146 5488 4558
rect 5552 4146 5580 5850
rect 5644 4622 5672 6394
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 5098 5764 6258
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5234 5856 5714
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 6012 4842 6040 7890
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5030 6132 5578
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5920 4814 6040 4842
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5828 4146 5856 4694
rect 5920 4622 5948 4814
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5368 3890 5396 4014
rect 5448 4004 5500 4010
rect 5632 4004 5684 4010
rect 5500 3964 5632 3992
rect 5448 3946 5500 3952
rect 5632 3946 5684 3952
rect 6012 3942 6040 4626
rect 5724 3936 5776 3942
rect 5368 3884 5724 3890
rect 6000 3936 6052 3942
rect 5368 3878 5776 3884
rect 5906 3904 5962 3913
rect 5368 3862 5764 3878
rect 5538 3768 5594 3777
rect 5538 3703 5594 3712
rect 5552 3670 5580 3703
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5552 3058 5580 3606
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5644 2854 5672 3862
rect 6000 3878 6052 3884
rect 5906 3839 5962 3848
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5000 2746 5120 2774
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 4252 1284 4304 1290
rect 4252 1226 4304 1232
rect 4264 800 4292 1226
rect 4632 800 4660 2042
rect 5000 800 5028 2746
rect 5736 2650 5764 3402
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5540 2644 5592 2650
rect 5724 2644 5776 2650
rect 5592 2604 5672 2632
rect 5540 2586 5592 2592
rect 5644 2530 5672 2604
rect 5724 2586 5776 2592
rect 5644 2502 5764 2530
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 2106 5212 2382
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5356 1556 5408 1562
rect 5356 1498 5408 1504
rect 5368 800 5396 1498
rect 5736 800 5764 2502
rect 5828 2446 5856 2790
rect 5920 2774 5948 3839
rect 6104 3058 6132 4966
rect 6196 3777 6224 9454
rect 6288 8974 6316 9522
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6182 3768 6238 3777
rect 6182 3703 6238 3712
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6288 2774 6316 8502
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6380 7410 6408 8026
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 5030 6408 7142
rect 6472 6390 6500 9386
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6564 8566 6592 8842
rect 6656 8634 6684 9522
rect 6748 9042 6776 10406
rect 7024 10266 7052 10610
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7116 10130 7144 10542
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6564 7818 6592 8502
rect 6840 8498 6868 8910
rect 6932 8634 6960 9930
rect 7300 9178 7328 10610
rect 7668 9586 7696 11222
rect 8404 11150 8432 11614
rect 8864 11354 8892 11698
rect 9048 11694 9076 13262
rect 10244 12986 10272 13874
rect 10980 13530 11008 15302
rect 11348 14346 11376 15370
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11348 13938 11376 14282
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 11072 12850 11100 13670
rect 11348 13258 11376 13874
rect 11532 13326 11560 14758
rect 11716 13530 11744 16050
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11808 14006 11836 15574
rect 12176 15502 12204 16594
rect 12636 16590 12664 19110
rect 12820 18766 12848 20538
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12728 16114 12756 16526
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15502 12296 15846
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12176 15026 12204 15438
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 11900 14074 11928 14962
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11354 9076 11494
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9416 11150 9444 11630
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10062 8156 10610
rect 8404 10470 8432 11086
rect 9140 10810 9168 11086
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9600 10674 9628 11494
rect 9968 10810 9996 12174
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10060 11082 10088 12038
rect 10612 11694 10640 12038
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7760 9722 7788 9998
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7470 9072 7526 9081
rect 7470 9007 7526 9016
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6918 8528 6974 8537
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6828 8492 6880 8498
rect 6918 8463 6974 8472
rect 6828 8434 6880 8440
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6472 5234 6500 6054
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6380 4593 6408 4694
rect 6366 4584 6422 4593
rect 6366 4519 6422 4528
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3126 6408 3878
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6564 2990 6592 6666
rect 6656 6497 6684 8434
rect 6840 7886 6868 8434
rect 6932 8294 6960 8463
rect 7024 8401 7052 8570
rect 7010 8392 7066 8401
rect 7010 8327 7066 8336
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 7342 6868 7482
rect 6932 7478 6960 7686
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6642 6488 6698 6497
rect 6642 6423 6698 6432
rect 6840 6118 6868 6598
rect 6932 6497 6960 7278
rect 7024 6984 7052 7346
rect 7104 6996 7156 7002
rect 7024 6956 7104 6984
rect 7104 6938 7156 6944
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6918 6488 6974 6497
rect 6918 6423 6974 6432
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6748 4146 6776 6054
rect 6932 5574 6960 6423
rect 7024 6322 7052 6598
rect 7208 6458 7236 6802
rect 7300 6730 7328 7686
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 7010 5536 7066 5545
rect 6932 5234 6960 5510
rect 7010 5471 7066 5480
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6748 3738 6776 4082
rect 6840 3942 6868 4558
rect 6932 4146 6960 4762
rect 7024 4214 7052 5471
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6748 3058 6776 3470
rect 7208 3210 7236 5578
rect 7392 5302 7420 8298
rect 7484 5545 7512 9007
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7470 5536 7526 5545
rect 7470 5471 7526 5480
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7392 4146 7420 4218
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 3398 7328 3674
rect 7392 3602 7420 4082
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 6828 3188 6880 3194
rect 7208 3182 7328 3210
rect 6828 3130 6880 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 5920 2746 6132 2774
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6104 800 6132 2746
rect 6196 2746 6316 2774
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6196 762 6224 2746
rect 6840 2650 6868 3130
rect 7196 3120 7248 3126
rect 7194 3088 7196 3097
rect 7248 3088 7250 3097
rect 7194 3023 7250 3032
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 6840 800 6868 2450
rect 7300 2378 7328 3182
rect 7392 2446 7420 3334
rect 7484 3097 7512 5170
rect 7576 4826 7604 8434
rect 7668 6254 7696 9522
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7760 9178 7788 9454
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 6798 7788 8910
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8514 8064 8774
rect 8404 8566 8432 10406
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8588 9518 8616 9590
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8772 8906 8800 9522
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8392 8560 8444 8566
rect 8036 8498 8156 8514
rect 8392 8502 8444 8508
rect 8036 8492 8168 8498
rect 8036 8486 8116 8492
rect 8116 8434 8168 8440
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 8090 7880 8298
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 8090 7972 8230
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7852 7886 7880 8026
rect 8956 7970 8984 10610
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9382 9076 9862
rect 9508 9722 9536 9930
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9036 8968 9088 8974
rect 9140 8956 9168 9386
rect 9088 8928 9168 8956
rect 9036 8910 9088 8916
rect 9048 8294 9076 8910
rect 9324 8673 9352 9590
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9042 9444 9454
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9310 8664 9366 8673
rect 9310 8599 9366 8608
rect 9508 8362 9536 9658
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 8956 7942 9168 7970
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7838 7576 7894 7585
rect 7838 7511 7894 7520
rect 7852 7478 7880 7511
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8116 7200 8168 7206
rect 8036 7160 8116 7188
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6254 7788 6734
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 6458 7880 6666
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7932 6316 7984 6322
rect 8036 6304 8064 7160
rect 8312 7177 8340 7210
rect 8116 7142 8168 7148
rect 8298 7168 8354 7177
rect 8298 7103 8354 7112
rect 8404 6458 8432 7754
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 7984 6276 8064 6304
rect 8116 6316 8168 6322
rect 7932 6258 7984 6264
rect 8116 6258 8168 6264
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 8128 5522 8156 6258
rect 8392 6248 8444 6254
rect 8390 6216 8392 6225
rect 8444 6216 8446 6225
rect 8390 6151 8446 6160
rect 8298 6080 8354 6089
rect 8298 6015 8354 6024
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 7944 5494 8156 5522
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7944 4622 7972 5494
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 8036 4282 8064 4490
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7576 4146 8064 4162
rect 7576 4140 8076 4146
rect 7576 4134 8024 4140
rect 7576 4078 7604 4134
rect 8024 4082 8076 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7840 4072 7892 4078
rect 8128 4026 8156 5306
rect 8220 4078 8248 5578
rect 8312 5098 8340 6015
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 7892 4020 8156 4026
rect 7840 4014 8156 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7852 3998 8156 4014
rect 7932 3936 7984 3942
rect 7984 3896 8156 3924
rect 7932 3878 7984 3884
rect 8128 3670 8156 3896
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7852 3346 7880 3470
rect 7852 3318 8064 3346
rect 8036 3194 8064 3318
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7470 3088 7526 3097
rect 7470 3023 7526 3032
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7196 1828 7248 1834
rect 7196 1770 7248 1776
rect 7208 800 7236 1770
rect 7576 800 7604 2994
rect 8128 2854 8156 3470
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 7944 800 7972 1362
rect 8312 800 8340 3839
rect 8390 3632 8446 3641
rect 8390 3567 8446 3576
rect 6196 734 6408 762
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8404 762 8432 3567
rect 8496 3194 8524 7346
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 5846 8708 6666
rect 8668 5840 8720 5846
rect 8666 5808 8668 5817
rect 8720 5808 8722 5817
rect 8666 5743 8722 5752
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8588 4214 8616 4694
rect 8680 4554 8708 5238
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 4282 8708 4490
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3602 8616 3878
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8574 3224 8630 3233
rect 8484 3188 8536 3194
rect 8574 3159 8576 3168
rect 8484 3130 8536 3136
rect 8628 3159 8630 3168
rect 8576 3130 8628 3136
rect 8680 3074 8708 4218
rect 8864 3602 8892 6938
rect 8956 6497 8984 7822
rect 9140 7750 9168 7942
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8942 6488 8998 6497
rect 8942 6423 8998 6432
rect 8956 6322 8984 6423
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8956 5846 8984 6122
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9048 5370 9076 7142
rect 9140 5710 9168 7686
rect 9324 7410 9352 8230
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6798 9352 7142
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9508 5574 9536 6831
rect 9600 6798 9628 10610
rect 9784 10266 9812 10610
rect 10612 10606 10640 11630
rect 10980 11082 11008 12650
rect 11348 12442 11376 13194
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11440 11898 11468 12718
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11624 11150 11652 12718
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9956 8968 10008 8974
rect 10048 8968 10100 8974
rect 9956 8910 10008 8916
rect 10046 8936 10048 8945
rect 10324 8968 10376 8974
rect 10100 8936 10102 8945
rect 9968 8634 9996 8910
rect 10324 8910 10376 8916
rect 10046 8871 10102 8880
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10336 8498 10364 8910
rect 10414 8800 10470 8809
rect 10414 8735 10470 8744
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9678 7848 9734 7857
rect 9678 7783 9734 7792
rect 9692 7002 9720 7783
rect 9784 7410 9812 8026
rect 10152 7528 10180 8434
rect 9876 7500 10180 7528
rect 10232 7540 10284 7546
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9770 7304 9826 7313
rect 9770 7239 9826 7248
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9692 6440 9720 6802
rect 9600 6412 9720 6440
rect 9600 6322 9628 6412
rect 9678 6352 9734 6361
rect 9588 6316 9640 6322
rect 9678 6287 9680 6296
rect 9588 6258 9640 6264
rect 9732 6287 9734 6296
rect 9680 6258 9732 6264
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9784 5302 9812 7239
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4826 9352 5170
rect 9770 4992 9826 5001
rect 9770 4927 9826 4936
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9784 4758 9812 4927
rect 9772 4752 9824 4758
rect 9876 4729 9904 7500
rect 10232 7482 10284 7488
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 6866 9996 7142
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10060 6338 10088 7278
rect 9968 6310 10088 6338
rect 9968 4978 9996 6310
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5166 10088 5510
rect 10152 5370 10180 7346
rect 10244 7274 10272 7482
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5710 10272 6258
rect 10336 6225 10364 6666
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10230 5536 10286 5545
rect 10230 5471 10286 5480
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9968 4950 10180 4978
rect 9772 4694 9824 4700
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8942 4176 8998 4185
rect 8942 4111 8998 4120
rect 8956 3942 8984 4111
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8944 3664 8996 3670
rect 9232 3652 9260 4558
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9588 4208 9640 4214
rect 9680 4208 9732 4214
rect 9588 4150 9640 4156
rect 9678 4176 9680 4185
rect 9732 4176 9734 4185
rect 9600 4060 9628 4150
rect 9678 4111 9734 4120
rect 9968 4078 9996 4490
rect 9956 4072 10008 4078
rect 9600 4032 9720 4060
rect 8996 3624 9260 3652
rect 8944 3606 8996 3612
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8496 3046 8708 3074
rect 8864 3058 8892 3538
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8852 3052 8904 3058
rect 8496 2378 8524 3046
rect 8852 2994 8904 3000
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8588 2446 8616 2790
rect 9048 2650 9076 3402
rect 9126 3088 9182 3097
rect 9126 3023 9128 3032
rect 9180 3023 9182 3032
rect 9128 2994 9180 3000
rect 9232 2854 9260 3624
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9324 2961 9352 3402
rect 9692 3398 9720 4032
rect 9956 4014 10008 4020
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9600 3058 9628 3334
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9496 2984 9548 2990
rect 9310 2952 9366 2961
rect 9968 2938 9996 4014
rect 10152 3346 10180 4950
rect 9548 2932 9996 2938
rect 9496 2926 9996 2932
rect 9508 2910 9996 2926
rect 9310 2887 9366 2896
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9416 2514 9444 2790
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9968 2446 9996 2910
rect 10060 3318 10180 3346
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9036 1148 9088 1154
rect 9036 1090 9088 1096
rect 8588 870 8708 898
rect 8588 762 8616 870
rect 8680 800 8708 870
rect 9048 800 9076 1090
rect 9416 800 9444 1974
rect 9784 870 9904 898
rect 9784 800 9812 870
rect 8404 734 8616 762
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 9876 762 9904 870
rect 10060 762 10088 3318
rect 10244 2774 10272 5471
rect 10336 5370 10364 6054
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10428 4865 10456 8735
rect 10612 7342 10640 10542
rect 10704 10062 10732 10950
rect 11808 10810 11836 12242
rect 11992 12238 12020 13262
rect 12176 12850 12204 14962
rect 12912 14346 12940 17206
rect 13004 16590 13032 17274
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13188 16522 13216 22066
rect 13372 22030 13400 23054
rect 13452 23044 13504 23050
rect 13452 22986 13504 22992
rect 13464 22438 13492 22986
rect 14844 22778 14872 23122
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 14292 21962 14320 22510
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14476 22098 14504 22374
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 20942 13492 21830
rect 13820 21480 13872 21486
rect 13740 21440 13820 21468
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13464 19446 13492 20470
rect 13740 20466 13768 21440
rect 13820 21422 13872 21428
rect 14292 21350 14320 21898
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13924 20058 13952 20402
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13464 18970 13492 19382
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13096 16250 13124 16458
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14618 13124 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 13188 14074 13216 14962
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13280 13938 13308 14214
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13372 13462 13400 18634
rect 13740 18290 13768 18702
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 16794 13768 17546
rect 13832 17338 13860 18634
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13832 16794 13860 17138
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 14016 16590 14044 17138
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16182 13492 16390
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13556 15994 13584 16118
rect 13464 15966 13584 15994
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13464 15162 13492 15966
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15706 13584 15846
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13464 14346 13492 15098
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12452 12442 12480 12854
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12636 12238 12664 13126
rect 13004 12986 13032 13194
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12434 13032 12582
rect 13004 12406 13124 12434
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10130 11100 10474
rect 11152 10464 11204 10470
rect 11204 10412 11376 10418
rect 11152 10406 11376 10412
rect 11164 10390 11376 10406
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10520 6118 10548 6666
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10414 4856 10470 4865
rect 10414 4791 10470 4800
rect 10520 4758 10548 6054
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10152 2746 10272 2774
rect 10152 800 10180 2746
rect 10336 1714 10364 3334
rect 10428 2650 10456 4150
rect 10612 3641 10640 6938
rect 10704 6866 10732 9998
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10784 9648 10836 9654
rect 10782 9616 10784 9625
rect 10836 9616 10838 9625
rect 11072 9586 11100 9930
rect 10782 9551 10838 9560
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10520 1902 10548 2382
rect 10704 2258 10732 6326
rect 10796 2922 10824 6938
rect 10888 5681 10916 8774
rect 10980 7750 11008 9386
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8498 11192 10390
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11256 10130 11284 10202
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 8566 11284 10066
rect 11348 10062 11376 10390
rect 11716 10266 11744 10610
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 8424 11112 8430
rect 11112 8372 11376 8378
rect 11060 8366 11376 8372
rect 11072 8350 11376 8366
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 6390 11008 7686
rect 11072 7410 11100 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11164 7410 11192 8026
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11256 6798 11284 7686
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5914 11008 6190
rect 11164 6186 11192 6598
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10874 5672 10930 5681
rect 10874 5607 10930 5616
rect 10966 5536 11022 5545
rect 10966 5471 11022 5480
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10796 2774 10824 2858
rect 10888 2836 10916 5238
rect 10980 5166 11008 5471
rect 11152 5228 11204 5234
rect 11072 5188 11152 5216
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10966 4856 11022 4865
rect 10966 4791 11022 4800
rect 10980 4758 11008 4791
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11072 4321 11100 5188
rect 11152 5170 11204 5176
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11058 4312 11114 4321
rect 11058 4247 11114 4256
rect 11164 3942 11192 4422
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11256 3534 11284 6394
rect 11348 5914 11376 8350
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11334 5400 11390 5409
rect 11334 5335 11390 5344
rect 11348 3942 11376 5335
rect 11440 5234 11468 9930
rect 11624 9586 11652 9930
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 8968 11572 8974
rect 11796 8968 11848 8974
rect 11572 8928 11744 8956
rect 11520 8910 11572 8916
rect 11716 8566 11744 8928
rect 11796 8910 11848 8916
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11612 8492 11664 8498
rect 11808 8480 11836 8910
rect 11900 8838 11928 11698
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12084 10062 12112 10202
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9926 12112 9998
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11992 8838 12020 9046
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12084 8548 12112 9862
rect 12268 9518 12296 11698
rect 12452 10606 12480 12106
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11762 13032 12038
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10062 12480 10542
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12268 9042 12296 9454
rect 12360 9110 12388 9590
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12452 8974 12480 9998
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12530 8800 12586 8809
rect 12530 8735 12586 8744
rect 11992 8520 12112 8548
rect 11888 8492 11940 8498
rect 11808 8452 11888 8480
rect 11612 8434 11664 8440
rect 11888 8434 11940 8440
rect 11532 7750 11560 8434
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11624 7546 11652 8434
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 7546 11928 7686
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11518 7440 11574 7449
rect 11518 7375 11574 7384
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11426 5128 11482 5137
rect 11426 5063 11482 5072
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10888 2808 11008 2836
rect 10796 2746 10916 2774
rect 10888 2378 10916 2746
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10704 2230 10916 2258
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10336 1686 10548 1714
rect 10520 800 10548 1686
rect 10888 800 10916 2230
rect 9876 734 10088 762
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 10980 762 11008 2808
rect 11440 2774 11468 5063
rect 11532 4321 11560 7375
rect 11992 6458 12020 8520
rect 12544 8362 12572 8735
rect 12636 8634 12664 11222
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12820 9586 12848 9930
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 8106 12480 8230
rect 12268 8078 12480 8106
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12084 7206 12112 7414
rect 12268 7410 12296 8078
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12544 7342 12572 7822
rect 12164 7336 12216 7342
rect 12532 7336 12584 7342
rect 12216 7284 12480 7290
rect 12164 7278 12480 7284
rect 12532 7278 12584 7284
rect 12176 7262 12480 7278
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12452 7002 12480 7262
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4826 11652 5170
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11518 4312 11574 4321
rect 11518 4247 11574 4256
rect 11624 4078 11652 4558
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11716 4146 11744 4218
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11532 2990 11560 3402
rect 11624 3058 11652 4014
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11808 2854 11836 6054
rect 11900 4282 11928 6287
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11992 5370 12020 5850
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4457 12020 4558
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 11978 4312 12034 4321
rect 11888 4276 11940 4282
rect 11978 4247 11980 4256
rect 11888 4218 11940 4224
rect 12032 4247 12034 4256
rect 11980 4218 12032 4224
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11888 3936 11940 3942
rect 11992 3913 12020 3946
rect 11888 3878 11940 3884
rect 11978 3904 12034 3913
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11900 2774 11928 3878
rect 11978 3839 12034 3848
rect 12084 3670 12112 6666
rect 12360 5914 12388 6938
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11980 3052 12032 3058
rect 12084 3040 12112 3606
rect 12032 3012 12112 3040
rect 11980 2994 12032 3000
rect 12176 2922 12204 4694
rect 12268 4486 12296 4694
rect 12360 4554 12388 5850
rect 12544 5778 12572 7278
rect 12636 6866 12664 8570
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12622 6352 12678 6361
rect 12622 6287 12624 6296
rect 12676 6287 12678 6296
rect 12624 6258 12676 6264
rect 12728 6254 12756 8502
rect 12820 8498 12848 9046
rect 12912 8838 12940 10542
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8838 13032 8910
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 7750 12940 8298
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 6798 12940 7686
rect 13096 6798 13124 12406
rect 13266 9616 13322 9625
rect 13372 9602 13400 13398
rect 13648 13326 13676 15982
rect 13636 13320 13688 13326
rect 14004 13320 14056 13326
rect 13636 13262 13688 13268
rect 14002 13288 14004 13297
rect 14056 13288 14058 13297
rect 14002 13223 14058 13232
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11150 13768 12242
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10606 13768 11086
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 9722 13768 10542
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13322 9574 13400 9602
rect 13266 9551 13322 9560
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13188 8906 13216 9046
rect 13176 8900 13228 8906
rect 13228 8860 13308 8888
rect 13176 8842 13228 8848
rect 13280 7206 13308 8860
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12820 6458 12848 6666
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 13096 6254 13124 6598
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12544 5234 12572 5714
rect 12636 5545 12664 6122
rect 12622 5536 12678 5545
rect 12622 5471 12678 5480
rect 12532 5228 12584 5234
rect 12452 5188 12532 5216
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12254 3768 12310 3777
rect 12254 3703 12256 3712
rect 12308 3703 12310 3712
rect 12256 3674 12308 3680
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 11440 2746 11652 2774
rect 11900 2746 12020 2774
rect 11164 870 11284 898
rect 11164 762 11192 870
rect 11256 800 11284 870
rect 11624 800 11652 2746
rect 11992 800 12020 2746
rect 12268 2582 12296 2926
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 2038 12296 2246
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12360 800 12388 3567
rect 12452 3534 12480 5188
rect 12532 5170 12584 5176
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12544 3534 12572 5034
rect 13096 4758 13124 5170
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4214 12848 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12714 4040 12770 4049
rect 12714 3975 12770 3984
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12452 3058 12480 3470
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12728 800 12756 3975
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 2446 13032 3470
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13096 800 13124 4218
rect 13188 4146 13216 6938
rect 13280 6662 13308 7142
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13372 6474 13400 9454
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13464 9081 13492 9114
rect 13450 9072 13506 9081
rect 13450 9007 13506 9016
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8566 13676 8910
rect 13740 8838 13768 9318
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13280 6458 13400 6474
rect 13268 6452 13400 6458
rect 13320 6446 13400 6452
rect 13268 6394 13320 6400
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13372 5710 13400 6326
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13464 4622 13492 6870
rect 13556 6662 13584 8434
rect 13648 7313 13676 8502
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13648 6798 13676 7239
rect 13740 6934 13768 8774
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5574 13676 6258
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13280 3738 13308 4150
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13280 3534 13308 3674
rect 13268 3528 13320 3534
rect 13174 3496 13230 3505
rect 13268 3470 13320 3476
rect 13174 3431 13176 3440
rect 13228 3431 13230 3440
rect 13176 3402 13228 3408
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13280 2106 13308 2246
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13556 800 13584 5306
rect 13832 2774 13860 13126
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12434 14044 12922
rect 13924 12406 14044 12434
rect 13924 10266 13952 12406
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 10810 14044 12174
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14108 10130 14136 19790
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 11898 14228 16594
rect 14292 15978 14320 21286
rect 14844 21146 14872 21490
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17338 14504 18022
rect 14568 17882 14596 18226
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14556 17672 14608 17678
rect 14740 17672 14792 17678
rect 14608 17620 14688 17626
rect 14556 17614 14688 17620
rect 14740 17614 14792 17620
rect 14936 17626 14964 25842
rect 15028 24614 15056 26318
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 15304 25362 15332 26182
rect 15488 25838 15516 27474
rect 15764 27470 15792 28562
rect 15948 28218 15976 29106
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 16132 28558 16160 28902
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 16868 28218 16896 29106
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15764 27062 15792 27406
rect 16868 27130 16896 28018
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15672 25838 15700 26250
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 15028 24274 15056 24550
rect 15212 24342 15240 24822
rect 15304 24750 15332 25298
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15108 21956 15160 21962
rect 15108 21898 15160 21904
rect 15120 21622 15148 21898
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15120 21010 15148 21558
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15120 20602 15148 20946
rect 15212 20942 15240 22374
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15304 21690 15332 21966
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15396 19922 15424 21830
rect 15488 21434 15516 25774
rect 15672 25242 15700 25774
rect 15764 25362 15792 26998
rect 17052 26994 17080 27474
rect 17420 27062 17448 29446
rect 17604 28014 17632 29582
rect 17788 29306 17816 29582
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 17972 28626 18000 29038
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 17868 28484 17920 28490
rect 17868 28426 17920 28432
rect 17880 28218 17908 28426
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17592 28008 17644 28014
rect 17592 27950 17644 27956
rect 17972 27946 18000 28562
rect 18064 28218 18092 29106
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18432 28994 18460 29038
rect 18524 29034 18552 29990
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 18248 28966 18460 28994
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18144 28552 18196 28558
rect 18248 28540 18276 28966
rect 18196 28512 18276 28540
rect 18144 28494 18196 28500
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 18156 28098 18184 28494
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18248 28150 18276 28358
rect 18064 28070 18184 28098
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 15948 26586 15976 26726
rect 15936 26580 15988 26586
rect 15936 26522 15988 26528
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15948 25974 15976 26318
rect 15936 25968 15988 25974
rect 15936 25910 15988 25916
rect 15752 25356 15804 25362
rect 15752 25298 15804 25304
rect 15672 25214 15792 25242
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15580 22030 15608 23598
rect 15672 23254 15700 23666
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 15672 22710 15700 23190
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15764 22642 15792 25214
rect 16040 24342 16068 26726
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15764 21554 15792 22578
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15488 21406 15608 21434
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 21146 15516 21286
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15580 21026 15608 21406
rect 15488 20998 15608 21026
rect 15488 20398 15516 20998
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15488 19802 15516 20334
rect 15580 20262 15608 20878
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19854 15608 20198
rect 15396 19774 15516 19802
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15396 19378 15424 19774
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15028 17746 15056 18362
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15120 17678 15148 19178
rect 15108 17672 15160 17678
rect 14568 17598 14688 17614
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14384 16590 14412 17206
rect 14568 17202 14596 17478
rect 14660 17218 14688 17598
rect 14752 17338 14780 17614
rect 14936 17598 15056 17626
rect 15108 17614 15160 17620
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14832 17264 14884 17270
rect 14660 17212 14832 17218
rect 14660 17206 14884 17212
rect 14556 17196 14608 17202
rect 14660 17190 14872 17206
rect 15028 17202 15056 17598
rect 15016 17196 15068 17202
rect 14556 17138 14608 17144
rect 15016 17138 15068 17144
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14384 16046 14412 16526
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14384 15570 14412 15982
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14476 15502 14504 16050
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14414 14412 14894
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14568 14056 14596 16118
rect 14476 14028 14596 14056
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 12434 14320 13670
rect 14476 13326 14504 14028
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 12986 14504 13262
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14292 12406 14412 12434
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9178 13952 9998
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14108 9024 14136 10066
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14292 9178 14320 9590
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14016 8996 14136 9024
rect 14016 8430 14044 8996
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 7410 14044 8230
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 6866 13952 7142
rect 13912 6860 13964 6866
rect 14108 6848 14136 8298
rect 14292 7970 14320 8366
rect 14200 7942 14320 7970
rect 14200 7206 14228 7942
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7546 14320 7822
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14384 7342 14412 12406
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14476 9450 14504 9522
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7886 14504 8230
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 13912 6802 13964 6808
rect 14016 6820 14136 6848
rect 14016 6390 14044 6820
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14108 5370 14136 6666
rect 14200 5846 14228 6666
rect 14188 5840 14240 5846
rect 14240 5800 14320 5828
rect 14188 5782 14240 5788
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13924 4060 13952 5102
rect 14108 4690 14136 5306
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14200 4185 14228 5578
rect 14292 4690 14320 5800
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4282 14320 4422
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14186 4176 14242 4185
rect 14292 4146 14320 4218
rect 14186 4111 14188 4120
rect 14240 4111 14242 4120
rect 14280 4140 14332 4146
rect 14188 4082 14240 4088
rect 14280 4082 14332 4088
rect 13924 4032 14044 4060
rect 13832 2746 13952 2774
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13832 2514 13860 2586
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13924 800 13952 2746
rect 10980 734 11192 762
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14016 762 14044 4032
rect 14292 4026 14320 4082
rect 14108 3998 14320 4026
rect 14108 3534 14136 3998
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3641 14320 3878
rect 14278 3632 14334 3641
rect 14278 3567 14334 3576
rect 14384 3534 14412 6938
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 2378 14136 3334
rect 14384 2922 14412 3470
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14476 2774 14504 7686
rect 14568 7546 14596 13874
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6322 14596 6598
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14660 5914 14688 17070
rect 14740 16584 14792 16590
rect 14936 16538 14964 17070
rect 15120 16998 15148 17614
rect 15396 17610 15424 19314
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18630 15516 18838
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15488 17066 15516 18566
rect 15580 18086 15608 19110
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17678 15792 18022
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14792 16532 14964 16538
rect 14740 16526 14964 16532
rect 14752 16510 14964 16526
rect 14844 16046 14872 16510
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14752 13682 14780 15982
rect 14844 15638 14872 15982
rect 15120 15978 15148 16934
rect 15764 16726 15792 17138
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15764 16590 15792 16662
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15672 16250 15700 16526
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14936 14074 14964 14962
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15212 13938 15240 15302
rect 15304 14346 15332 15846
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15396 13870 15424 14826
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 14752 13654 14872 13682
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 12918 14780 13126
rect 14844 12986 14872 13654
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14844 12238 14872 12922
rect 14936 12442 14964 13262
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 12889 15424 13126
rect 15382 12880 15438 12889
rect 15382 12815 15438 12824
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15028 11082 15056 12106
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15120 11121 15148 11834
rect 15212 11150 15240 11834
rect 15304 11762 15332 12582
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15488 11354 15516 12786
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15580 11150 15608 12174
rect 15672 11694 15700 14214
rect 15764 13870 15792 15846
rect 15856 15502 15884 23802
rect 16224 23730 16252 26930
rect 16868 26586 16896 26930
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 16224 22030 16252 23122
rect 16316 22642 16344 25298
rect 16868 24410 16896 25842
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16316 22522 16344 22578
rect 16316 22494 16436 22522
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21622 16344 21830
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16408 21418 16436 22494
rect 16500 21894 16528 24142
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16592 23254 16620 24074
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16684 23322 16712 23462
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16776 23066 16804 23802
rect 16960 23662 16988 24142
rect 17052 24138 17080 26930
rect 17420 26314 17448 26998
rect 17512 26314 17540 27406
rect 17972 27062 18000 27882
rect 18064 27470 18092 28070
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18156 27606 18184 27950
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 18340 26586 18368 27950
rect 18800 27878 18828 28426
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17500 26308 17552 26314
rect 17500 26250 17552 26256
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17236 24954 17264 25094
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16684 23038 16804 23066
rect 16684 22506 16712 23038
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21690 16528 21830
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16408 21146 16436 21354
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18290 15976 18634
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16040 17202 16068 20810
rect 16408 20466 16436 21082
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16592 20942 16620 21014
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16224 18290 16252 19790
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16408 18970 16436 19722
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16592 18766 16620 19110
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 17610 16252 18226
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 15570 15976 16050
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15200 11144 15252 11150
rect 15106 11112 15162 11121
rect 15016 11076 15068 11082
rect 15200 11086 15252 11092
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15106 11047 15162 11056
rect 15016 11018 15068 11024
rect 15028 10742 15056 11018
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15120 10674 15148 11047
rect 15580 10674 15608 11086
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15120 9926 15148 10202
rect 15580 10130 15608 10610
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15212 9518 15240 9590
rect 15200 9512 15252 9518
rect 15252 9472 15332 9500
rect 15200 9454 15252 9460
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14568 4826 14596 5578
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14568 4010 14596 4762
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4214 14688 4422
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14646 4040 14702 4049
rect 14556 4004 14608 4010
rect 14646 3975 14702 3984
rect 14556 3946 14608 3952
rect 14568 3602 14596 3946
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14660 3534 14688 3975
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14476 2746 14688 2774
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14200 870 14320 898
rect 14200 762 14228 870
rect 14292 800 14320 870
rect 14660 800 14688 2746
rect 14016 734 14228 762
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 14752 762 14780 7482
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14844 7274 14872 7346
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14936 7154 14964 9318
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15028 7410 15056 7822
rect 15212 7546 15240 8434
rect 15304 7954 15332 9472
rect 15396 8945 15424 9998
rect 15672 9586 15700 10950
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15764 9024 15792 12786
rect 15488 8996 15792 9024
rect 15382 8936 15438 8945
rect 15382 8871 15438 8880
rect 15396 8430 15424 8871
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15396 8022 15424 8366
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15028 7313 15056 7346
rect 15014 7304 15070 7313
rect 15014 7239 15070 7248
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 14844 7126 14964 7154
rect 14844 6118 14872 7126
rect 15120 6390 15148 7210
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15016 6316 15068 6322
rect 14936 6276 15016 6304
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14936 5846 14964 6276
rect 15016 6258 15068 6264
rect 15016 6112 15068 6118
rect 15212 6066 15240 7346
rect 15382 6896 15438 6905
rect 15382 6831 15438 6840
rect 15396 6458 15424 6831
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6338 15516 8996
rect 15856 8922 15884 13262
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15580 8894 15884 8922
rect 15580 7750 15608 8894
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15672 7478 15700 8774
rect 15948 7970 15976 13126
rect 16040 12442 16068 17138
rect 16224 17066 16252 17546
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 14618 16160 15982
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16224 14414 16252 17002
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16408 15502 16436 15574
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 12714 16252 14350
rect 16408 14006 16436 15438
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16040 11150 16068 12378
rect 16224 12306 16252 12650
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16132 11082 16160 12106
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15764 7942 15976 7970
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15764 7324 15792 7942
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15566 7304 15622 7313
rect 15566 7239 15622 7248
rect 15672 7296 15792 7324
rect 15580 6390 15608 7239
rect 15016 6054 15068 6060
rect 15028 5914 15056 6054
rect 15120 6038 15240 6066
rect 15304 6310 15516 6338
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 15120 5778 15148 6038
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 4214 14964 5578
rect 15212 5234 15240 5850
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15120 4706 15148 5170
rect 15212 4826 15240 5170
rect 15304 5166 15332 6310
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 5302 15424 5646
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15120 4678 15240 4706
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14844 3466 14872 3567
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14936 3194 14964 4150
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15028 2514 15056 4490
rect 15120 3602 15148 4558
rect 15212 4282 15240 4678
rect 15304 4622 15332 4966
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15292 4072 15344 4078
rect 15396 4060 15424 5102
rect 15476 5024 15528 5030
rect 15474 4992 15476 5001
rect 15528 4992 15530 5001
rect 15474 4927 15530 4936
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15344 4032 15424 4060
rect 15292 4014 15344 4020
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15212 2650 15240 3470
rect 15396 3466 15424 3674
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 14936 870 15056 898
rect 14936 762 14964 870
rect 15028 800 15056 870
rect 15396 800 15424 2994
rect 15580 2514 15608 4626
rect 15672 4010 15700 7296
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15764 6186 15792 6666
rect 15856 6458 15884 7346
rect 15948 7002 15976 7822
rect 16040 7546 16068 7958
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 6458 15976 6666
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15936 6452 15988 6458
rect 16132 6440 16160 10066
rect 16316 9602 16344 12038
rect 16500 11150 16528 15642
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16592 15366 16620 15574
rect 16684 15502 16712 22442
rect 16776 22098 16804 22918
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16960 21554 16988 23462
rect 17040 23180 17092 23186
rect 17144 23168 17172 24686
rect 17236 24138 17264 24890
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17092 23140 17172 23168
rect 17040 23122 17092 23128
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 17144 22234 17172 22510
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 19530 16804 20878
rect 16960 20398 16988 21014
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16960 19854 16988 20334
rect 17052 19922 17080 20878
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16776 19502 16896 19530
rect 16868 19378 16896 19502
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16776 17218 16804 19246
rect 16868 18630 16896 19314
rect 16960 18834 16988 19654
rect 17052 19378 17080 19858
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 17882 16896 18566
rect 17052 18222 17080 19314
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17052 17882 17080 18022
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16776 17190 16896 17218
rect 17144 17202 17172 19382
rect 17236 19378 17264 24074
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17328 21962 17356 22918
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 17328 21350 17356 21898
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17328 19990 17356 21286
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17236 18766 17264 19178
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17236 17678 17264 18702
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17542 17264 17614
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16776 16250 16804 17070
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16776 16114 16804 16186
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16776 15722 16804 16050
rect 16868 15881 16896 17190
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16960 16794 16988 17138
rect 17144 16998 17172 17138
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16854 15872 16910 15881
rect 16854 15807 16910 15816
rect 16776 15694 16896 15722
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 14074 16712 14282
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11150 16620 11494
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16684 11257 16712 11290
rect 16670 11248 16726 11257
rect 16670 11183 16726 11192
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16316 9574 16436 9602
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 8090 16252 8434
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16224 7886 16252 8026
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15936 6394 15988 6400
rect 16040 6412 16160 6440
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15764 800 15792 5782
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15948 5234 15976 5578
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15856 3126 15884 3538
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 16040 3058 16068 6412
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16132 5914 16160 6258
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16120 5772 16172 5778
rect 16224 5760 16252 6598
rect 16302 6216 16358 6225
rect 16302 6151 16358 6160
rect 16172 5732 16252 5760
rect 16120 5714 16172 5720
rect 16316 4282 16344 6151
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 15948 2310 15976 2586
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 16132 800 16160 2790
rect 16224 2446 16252 4014
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16408 2106 16436 9574
rect 16500 9518 16528 9998
rect 16592 9722 16620 10542
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16684 8362 16712 9658
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 5234 16528 7142
rect 16592 5710 16620 7414
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6118 16712 6598
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16776 5556 16804 15506
rect 16868 15450 16896 15694
rect 16960 15570 16988 16458
rect 17144 16454 17172 16594
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16868 15422 16988 15450
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 13938 16896 15302
rect 16960 15026 16988 15422
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 15026 17172 15370
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16960 12918 16988 14962
rect 17144 14482 17172 14962
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 11354 16896 12786
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 11014 16896 11086
rect 16856 11008 16908 11014
rect 16960 10985 16988 11698
rect 17052 11354 17080 12922
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17040 11008 17092 11014
rect 16856 10950 16908 10956
rect 16946 10976 17002 10985
rect 17040 10950 17092 10956
rect 16946 10911 17002 10920
rect 16960 10266 16988 10911
rect 17052 10674 17080 10950
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 9722 16896 9930
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 9217 16896 9522
rect 16960 9489 16988 10202
rect 16946 9480 17002 9489
rect 16946 9415 17002 9424
rect 16854 9208 16910 9217
rect 16854 9143 16910 9152
rect 16960 8974 16988 9415
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16960 8498 16988 8910
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17052 7834 17080 8910
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16960 7806 17080 7834
rect 16868 5778 16896 7754
rect 16960 5846 16988 7806
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17052 5574 17080 7686
rect 17040 5568 17092 5574
rect 16776 5528 16988 5556
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16684 4554 16712 4694
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16684 4185 16712 4490
rect 16670 4176 16726 4185
rect 16670 4111 16726 4120
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16684 2514 16712 3878
rect 16776 3777 16804 4490
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16868 3194 16896 4082
rect 16960 3738 16988 5528
rect 17040 5510 17092 5516
rect 17040 3936 17092 3942
rect 17038 3904 17040 3913
rect 17092 3904 17094 3913
rect 17038 3839 17094 3848
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17144 2774 17172 13738
rect 17236 13462 17264 17478
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17328 12434 17356 18770
rect 17420 16522 17448 26250
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17512 25294 17540 25638
rect 18052 25424 18104 25430
rect 18052 25366 18104 25372
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24206 17540 24550
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17604 22982 17632 23054
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17788 21690 17816 24142
rect 17880 23730 17908 24822
rect 17972 24750 18000 25094
rect 18064 24818 18092 25366
rect 18248 25294 18276 26318
rect 18604 26308 18656 26314
rect 18604 26250 18656 26256
rect 18616 25906 18644 26250
rect 18696 25968 18748 25974
rect 18696 25910 18748 25916
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18512 25832 18564 25838
rect 18564 25780 18644 25786
rect 18512 25774 18644 25780
rect 18524 25758 18644 25774
rect 18420 25696 18472 25702
rect 18420 25638 18472 25644
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 18248 24614 18276 25230
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18064 23322 18092 23666
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18052 23180 18104 23186
rect 18052 23122 18104 23128
rect 18064 22094 18092 23122
rect 18156 23118 18184 23666
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18248 22710 18276 24006
rect 18340 23186 18368 24278
rect 18432 23662 18460 25638
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18524 24070 18552 24754
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23730 18552 24006
rect 18616 23866 18644 25758
rect 18708 24954 18736 25910
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18420 23656 18472 23662
rect 18616 23610 18644 23802
rect 18420 23598 18472 23604
rect 18524 23582 18644 23610
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18340 22778 18368 22918
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18144 22094 18196 22098
rect 18524 22094 18552 23582
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22438 18644 22986
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18064 22092 18196 22094
rect 18064 22066 18144 22092
rect 18144 22034 18196 22040
rect 18248 22066 18552 22094
rect 18248 22030 18276 22066
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17696 19854 17724 20810
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18064 20534 18092 20742
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17696 18766 17724 19790
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17696 18630 17724 18702
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17788 17626 17816 19790
rect 17880 18834 17908 19858
rect 18156 19310 18184 21490
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18432 20618 18460 20878
rect 18432 20602 18552 20618
rect 18432 20596 18564 20602
rect 18432 20590 18512 20596
rect 18512 20538 18564 20544
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19378 18368 19654
rect 18524 19378 18552 20538
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17880 17746 17908 18770
rect 18524 18698 18552 19314
rect 18616 18766 18644 22374
rect 18800 22094 18828 27814
rect 19076 27130 19104 29106
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28098 19196 28970
rect 19260 28540 19288 29106
rect 19892 29096 19944 29102
rect 19892 29038 19944 29044
rect 19904 28558 19932 29038
rect 19996 28762 20024 29582
rect 20456 29170 20484 29990
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20456 29050 20484 29106
rect 20364 29022 20484 29050
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19340 28552 19392 28558
rect 19260 28512 19340 28540
rect 19260 28218 19288 28512
rect 19340 28494 19392 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19168 28082 19288 28098
rect 19168 28076 19300 28082
rect 19168 28070 19248 28076
rect 19248 28018 19300 28024
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19168 27470 19196 27950
rect 19156 27464 19208 27470
rect 19156 27406 19208 27412
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19168 27062 19196 27406
rect 19156 27056 19208 27062
rect 19156 26998 19208 27004
rect 19260 26874 19288 28018
rect 19444 27606 19472 28426
rect 19996 28393 20024 28426
rect 19982 28384 20038 28393
rect 19574 28316 19882 28336
rect 19982 28319 20038 28328
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 18984 26846 19288 26874
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18892 24274 18920 24686
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18708 22066 18828 22094
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17762 18000 18090
rect 18156 17882 18184 18294
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18524 17814 18552 18634
rect 18512 17808 18564 17814
rect 17868 17740 17920 17746
rect 17972 17734 18184 17762
rect 18512 17750 18564 17756
rect 17868 17682 17920 17688
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17512 15366 17540 17478
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17604 16454 17632 16526
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17512 14770 17540 15302
rect 17420 14742 17540 14770
rect 17420 13818 17448 14742
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17512 13938 17540 14554
rect 17604 14550 17632 16390
rect 17696 16114 17724 17614
rect 17788 17598 17908 17626
rect 17774 17504 17830 17513
rect 17774 17439 17830 17448
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17682 15872 17738 15881
rect 17682 15807 17738 15816
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17604 13938 17632 14486
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17420 13790 17632 13818
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17328 12406 17448 12434
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17224 9376 17276 9382
rect 17222 9344 17224 9353
rect 17276 9344 17278 9353
rect 17222 9279 17278 9288
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 6458 17264 7346
rect 17328 6610 17356 11290
rect 17420 10554 17448 12406
rect 17512 12238 17540 12582
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17604 11898 17632 13790
rect 17696 13734 17724 15807
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17512 11150 17540 11290
rect 17604 11150 17632 11494
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17420 10526 17632 10554
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 8566 17448 10406
rect 17498 9616 17554 9625
rect 17498 9551 17554 9560
rect 17512 9518 17540 9551
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 8906 17540 9318
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17604 8650 17632 10526
rect 17696 8974 17724 13398
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17604 8622 17724 8650
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17604 7886 17632 8502
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7478 17632 7822
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17590 6760 17646 6769
rect 17590 6695 17646 6704
rect 17328 6582 17540 6610
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17328 6338 17356 6394
rect 17236 6310 17356 6338
rect 17236 5778 17264 6310
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17236 5114 17264 5714
rect 17236 5086 17448 5114
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4146 17264 4966
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 3738 17356 4490
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17420 3398 17448 5086
rect 17512 4842 17540 6582
rect 17604 6322 17632 6695
rect 17696 6390 17724 8622
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17788 6202 17816 17439
rect 17880 16674 17908 17598
rect 17880 16646 18000 16674
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17880 16250 17908 16526
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17972 16182 18000 16646
rect 18156 16590 18184 17734
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18144 16584 18196 16590
rect 18196 16532 18276 16538
rect 18144 16526 18276 16532
rect 18156 16510 18276 16526
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 18248 16046 18276 16510
rect 18616 16114 18644 16594
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 15910 18276 15982
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17972 15094 18000 15506
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14482 17908 14894
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 14006 17908 14418
rect 17972 14414 18000 15030
rect 18156 15026 18184 15438
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 11558 17908 13670
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 11286 17908 11494
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10985 17908 11086
rect 17866 10976 17922 10985
rect 17866 10911 17922 10920
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 10130 17908 10542
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17880 7818 17908 10066
rect 17972 9586 18000 13806
rect 18064 12782 18092 14758
rect 18156 14278 18184 14962
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 13326 18184 14214
rect 18248 14074 18276 15846
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 14408 18472 14414
rect 18340 14368 18420 14396
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18248 12918 18276 13126
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 11830 18092 12038
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 7886 18000 9318
rect 18064 8634 18092 11630
rect 18248 10810 18276 12174
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18156 8090 18184 10610
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 8294 18276 9522
rect 18340 9042 18368 14368
rect 18420 14350 18472 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13326 18460 14214
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18524 11626 18552 15438
rect 18616 15094 18644 16050
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18616 14482 18644 15030
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18616 13988 18644 14418
rect 18708 14414 18736 22066
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18800 19378 18828 19722
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18800 17490 18828 19314
rect 18892 17678 18920 24210
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18800 17462 18920 17490
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18696 14000 18748 14006
rect 18616 13960 18696 13988
rect 18696 13942 18748 13948
rect 18694 13832 18750 13841
rect 18694 13767 18750 13776
rect 18708 13734 18736 13767
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18510 11248 18566 11257
rect 18510 11183 18566 11192
rect 18524 11150 18552 11183
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18432 10266 18460 11086
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18340 8809 18368 8842
rect 18326 8800 18382 8809
rect 18326 8735 18382 8744
rect 18432 8673 18460 9930
rect 18604 9580 18656 9586
rect 18524 9540 18604 9568
rect 18524 9178 18552 9540
rect 18604 9522 18656 9528
rect 18602 9208 18658 9217
rect 18512 9172 18564 9178
rect 18602 9143 18604 9152
rect 18512 9114 18564 9120
rect 18656 9143 18658 9152
rect 18604 9114 18656 9120
rect 18524 8974 18552 9114
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18708 8838 18736 11494
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18418 8664 18474 8673
rect 18418 8599 18474 8608
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17604 6174 17816 6202
rect 17604 5778 17632 6174
rect 17880 5794 17908 6666
rect 18064 6254 18092 6734
rect 18432 6730 18460 7414
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17696 5766 17908 5794
rect 17972 5778 18000 6054
rect 18064 5778 18092 6190
rect 17960 5772 18012 5778
rect 17696 5710 17724 5766
rect 17960 5714 18012 5720
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17972 5166 18000 5714
rect 18432 5710 18460 6666
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17512 4814 17632 4842
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 16868 2746 17172 2774
rect 17420 2774 17448 3334
rect 17420 2746 17540 2774
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16500 800 16528 2246
rect 16868 800 16896 2746
rect 17512 2582 17540 2746
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17236 800 17264 2518
rect 17604 800 17632 4814
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 2650 17724 4422
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18064 3126 18092 4218
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 18064 2446 18092 3062
rect 18156 2650 18184 4490
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3641 18276 4014
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18234 3632 18290 3641
rect 18234 3567 18236 3576
rect 18288 3567 18290 3576
rect 18236 3538 18288 3544
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18248 2854 18276 3402
rect 18340 2922 18368 3674
rect 18524 2972 18552 8502
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6390 18644 7142
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18616 3670 18644 4014
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18524 2944 18644 2972
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18340 2446 18368 2858
rect 18616 2650 18644 2944
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18616 2038 18644 2382
rect 18604 2032 18656 2038
rect 18604 1974 18656 1980
rect 18328 1760 18380 1766
rect 18328 1702 18380 1708
rect 17960 1420 18012 1426
rect 17960 1362 18012 1368
rect 17972 800 18000 1362
rect 18340 800 18368 1702
rect 18708 800 18736 4966
rect 18800 3738 18828 16526
rect 18892 13734 18920 17462
rect 18984 13938 19012 26846
rect 19352 26586 19380 27474
rect 19996 27334 20024 28319
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 19984 27328 20036 27334
rect 19982 27296 19984 27305
rect 20036 27296 20038 27305
rect 19574 27228 19882 27248
rect 19982 27231 20038 27240
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 20180 27130 20208 27950
rect 20272 27674 20300 28018
rect 20260 27668 20312 27674
rect 20260 27610 20312 27616
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19076 21146 19104 26386
rect 19260 24750 19288 26454
rect 19812 26382 19840 26998
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19800 26376 19852 26382
rect 20168 26376 20220 26382
rect 19852 26324 20024 26330
rect 19800 26318 20024 26324
rect 20168 26318 20220 26324
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19260 24154 19288 24686
rect 19352 24274 19380 26318
rect 19812 26302 20024 26318
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19904 25498 19932 25638
rect 19892 25492 19944 25498
rect 19892 25434 19944 25440
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19444 24206 19472 25230
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24818 20024 26302
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 20088 25906 20116 25978
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19890 24304 19946 24313
rect 19890 24239 19946 24248
rect 19904 24206 19932 24239
rect 20088 24206 20116 25842
rect 19432 24200 19484 24206
rect 19156 24132 19208 24138
rect 19260 24126 19380 24154
rect 19432 24142 19484 24148
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19156 24074 19208 24080
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19168 20942 19196 24074
rect 19352 23338 19380 24126
rect 19444 23508 19472 24142
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23798 20024 24006
rect 20088 23798 20116 24142
rect 20180 24070 20208 26318
rect 20272 25362 20300 26930
rect 20364 26858 20392 29022
rect 20352 26852 20404 26858
rect 20352 26794 20404 26800
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19524 23520 19576 23526
rect 19444 23480 19524 23508
rect 19524 23462 19576 23468
rect 19352 23310 19472 23338
rect 19444 23186 19472 23310
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19340 23112 19392 23118
rect 19260 23060 19340 23066
rect 19536 23066 19564 23462
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19628 23118 19656 23258
rect 19260 23054 19392 23060
rect 19260 23038 19380 23054
rect 19444 23038 19564 23066
rect 19616 23112 19668 23118
rect 19892 23112 19944 23118
rect 19616 23054 19668 23060
rect 19890 23080 19892 23089
rect 19944 23080 19946 23089
rect 19260 22710 19288 23038
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19352 22166 19380 22578
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19340 22024 19392 22030
rect 19444 22012 19472 23038
rect 19890 23015 19946 23024
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 22234 19564 22374
rect 19996 22234 20024 23598
rect 20088 22642 20116 23734
rect 20180 23730 20208 24006
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20074 22536 20130 22545
rect 20074 22471 20130 22480
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19392 21984 19472 22012
rect 19340 21966 19392 21972
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19076 20330 19104 20878
rect 19260 20618 19288 21286
rect 19352 21010 19380 21966
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21146 20024 21830
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 20088 20942 20116 22471
rect 20180 22166 20208 23122
rect 20272 22506 20300 25298
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20364 22386 20392 26794
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20456 23720 20484 26318
rect 20444 23714 20496 23720
rect 20444 23656 20496 23662
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20456 23322 20484 23530
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20272 22358 20392 22386
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 20180 21690 20208 22102
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19168 20590 19288 20618
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19168 19310 19196 20590
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19260 19446 19288 20402
rect 20272 19938 20300 22358
rect 20350 22264 20406 22273
rect 20350 22199 20406 22208
rect 20180 19910 20300 19938
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20074 19816 20130 19825
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19553 20024 19790
rect 20074 19751 20130 19760
rect 19982 19544 20038 19553
rect 19982 19479 20038 19488
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 20088 19378 20116 19751
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19904 18970 19932 19314
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19430 18864 19486 18873
rect 19430 18799 19486 18808
rect 19444 18766 19472 18799
rect 19432 18760 19484 18766
rect 19984 18760 20036 18766
rect 19432 18702 19484 18708
rect 19798 18728 19854 18737
rect 19340 18692 19392 18698
rect 19984 18702 20036 18708
rect 19798 18663 19800 18672
rect 19340 18634 19392 18640
rect 19852 18663 19854 18672
rect 19800 18634 19852 18640
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 19076 13802 19104 18158
rect 19260 17882 19288 18226
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16726 19196 17070
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19168 16250 19196 16458
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19260 15570 19288 16934
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19352 13977 19380 18634
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 17678 19472 18566
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18426 20024 18702
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19536 18193 19564 18294
rect 19522 18184 19578 18193
rect 19522 18119 19578 18128
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19536 17746 19564 18022
rect 19628 17785 19656 18022
rect 19614 17776 19670 17785
rect 19524 17740 19576 17746
rect 19614 17711 19670 17720
rect 19524 17682 19576 17688
rect 20088 17678 20116 19110
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19444 14890 19472 17206
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19536 16697 19564 17138
rect 19996 16794 20024 17138
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20088 16726 20116 17614
rect 20076 16720 20128 16726
rect 19522 16688 19578 16697
rect 20076 16662 20128 16668
rect 19522 16623 19578 16632
rect 19524 16584 19576 16590
rect 19522 16552 19524 16561
rect 19576 16552 19578 16561
rect 19522 16487 19578 16496
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 19616 16040 19668 16046
rect 19720 16017 19748 16118
rect 19892 16108 19944 16114
rect 20076 16108 20128 16114
rect 19944 16068 20024 16096
rect 19892 16050 19944 16056
rect 19616 15982 19668 15988
rect 19706 16008 19762 16017
rect 19628 15745 19656 15982
rect 19706 15943 19762 15952
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19614 15736 19670 15745
rect 19614 15671 19670 15680
rect 19812 15570 19840 15914
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19524 14952 19576 14958
rect 19522 14920 19524 14929
rect 19576 14920 19578 14929
rect 19432 14884 19484 14890
rect 19522 14855 19578 14864
rect 19892 14884 19944 14890
rect 19432 14826 19484 14832
rect 19892 14826 19944 14832
rect 19904 14657 19932 14826
rect 19890 14648 19946 14657
rect 19890 14583 19946 14592
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19338 13968 19394 13977
rect 19338 13903 19394 13912
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18880 13728 18932 13734
rect 19248 13728 19300 13734
rect 18880 13670 18932 13676
rect 19154 13696 19210 13705
rect 19248 13670 19300 13676
rect 19154 13631 19210 13640
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18892 9382 18920 9862
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18878 9072 18934 9081
rect 18878 9007 18880 9016
rect 18932 9007 18934 9016
rect 18880 8978 18932 8984
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18892 4146 18920 8298
rect 18984 5352 19012 11562
rect 19076 10198 19104 11698
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19064 9512 19116 9518
rect 19062 9480 19064 9489
rect 19116 9480 19118 9489
rect 19062 9415 19118 9424
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19076 8498 19104 8842
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19076 7818 19104 8434
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 18984 5324 19104 5352
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18984 3738 19012 5170
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19076 3466 19104 5324
rect 19168 4146 19196 13631
rect 19260 11694 19288 13670
rect 19444 13394 19472 14350
rect 19536 14260 19564 14486
rect 19996 14482 20024 16068
rect 20076 16050 20128 16056
rect 20088 14890 20116 16050
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19505 14232 19564 14260
rect 19505 14056 19533 14232
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19505 14028 19656 14056
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19536 13433 19564 13874
rect 19628 13734 19656 14028
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19996 13530 20024 14418
rect 20180 13938 20208 19910
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20272 19514 20300 19790
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20272 15638 20300 19246
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 14940 20300 15438
rect 20364 15094 20392 22199
rect 20456 21554 20484 23258
rect 20548 22030 20576 46514
rect 24872 35894 24900 46990
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 24872 35866 24992 35894
rect 20996 30728 21048 30734
rect 20996 30670 21048 30676
rect 21008 29850 21036 30670
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 20640 28762 20668 29650
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20824 29306 20852 29582
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20628 28756 20680 28762
rect 20628 28698 20680 28704
rect 20628 28416 20680 28422
rect 20628 28358 20680 28364
rect 20640 28218 20668 28358
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20824 28014 20852 28902
rect 21088 28484 21140 28490
rect 21088 28426 21140 28432
rect 21100 28218 21128 28426
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 21284 28082 21312 29446
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22664 28762 22692 29106
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 21824 28416 21876 28422
rect 21822 28384 21824 28393
rect 21876 28384 21878 28393
rect 21822 28319 21878 28328
rect 22112 28082 22140 28494
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21364 28076 21416 28082
rect 21364 28018 21416 28024
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20824 27334 20852 27950
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20640 24818 20668 25842
rect 20732 25838 20760 26930
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20720 25832 20772 25838
rect 20720 25774 20772 25780
rect 20732 25430 20760 25774
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20824 25294 20852 25842
rect 20916 25702 20944 26522
rect 21284 25922 21312 27270
rect 21376 26042 21404 28018
rect 21824 27872 21876 27878
rect 21824 27814 21876 27820
rect 21836 27538 21864 27814
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21652 26382 21680 26862
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21284 25894 21404 25922
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20916 25498 20944 25638
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 24410 20668 24550
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20732 23730 20760 25162
rect 20824 24818 20852 25230
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20824 24206 20852 24754
rect 20916 24682 20944 25434
rect 21284 25430 21312 25774
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 20904 24676 20956 24682
rect 20904 24618 20956 24624
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20732 23186 20760 23666
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20640 22710 20668 23054
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20640 21690 20668 21966
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20732 21554 20760 22374
rect 20444 21548 20496 21554
rect 20720 21548 20772 21554
rect 20444 21490 20496 21496
rect 20640 21508 20720 21536
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20456 16674 20484 20334
rect 20548 20058 20576 20742
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19854 20668 21508
rect 20720 21490 20772 21496
rect 20720 19984 20772 19990
rect 20718 19952 20720 19961
rect 20772 19952 20774 19961
rect 20718 19887 20774 19896
rect 20628 19848 20680 19854
rect 20824 19825 20852 24142
rect 21284 23730 21312 25366
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 22642 21036 23462
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20916 22098 20944 22578
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 20628 19790 20680 19796
rect 20810 19816 20866 19825
rect 20536 19372 20588 19378
rect 20640 19360 20668 19790
rect 20720 19780 20772 19786
rect 20810 19751 20866 19760
rect 20720 19722 20772 19728
rect 20588 19332 20668 19360
rect 20536 19314 20588 19320
rect 20548 17678 20576 19314
rect 20732 18902 20760 19722
rect 20916 19394 20944 22034
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 20534 21036 21286
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 21008 19514 21036 20470
rect 21100 20466 21128 22714
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21192 20398 21220 23122
rect 21284 22778 21312 23666
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22234 21312 22578
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21376 22114 21404 25894
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21560 24274 21588 24754
rect 21836 24410 21864 26794
rect 22020 26246 22048 28018
rect 22112 27538 22140 28018
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 21916 24744 21968 24750
rect 21968 24704 22048 24732
rect 21916 24686 21968 24692
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21284 22086 21404 22114
rect 21180 20392 21232 20398
rect 21100 20340 21180 20346
rect 21100 20334 21232 20340
rect 21100 20318 21220 20334
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20824 19378 20944 19394
rect 20812 19372 20944 19378
rect 20864 19366 20944 19372
rect 20996 19372 21048 19378
rect 20812 19314 20864 19320
rect 20996 19314 21048 19320
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20824 18766 20852 19314
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20628 18760 20680 18766
rect 20812 18760 20864 18766
rect 20628 18702 20680 18708
rect 20718 18728 20774 18737
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20640 17270 20668 18702
rect 20812 18702 20864 18708
rect 20718 18663 20774 18672
rect 20732 18154 20760 18663
rect 20824 18630 20852 18702
rect 20916 18698 20944 18906
rect 21008 18766 21036 19314
rect 21100 18834 21128 20318
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19718 21220 20198
rect 21284 20074 21312 22086
rect 21456 20868 21508 20874
rect 21456 20810 21508 20816
rect 21284 20046 21404 20074
rect 21468 20058 21496 20810
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21178 19544 21234 19553
rect 21178 19479 21234 19488
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 20996 18760 21048 18766
rect 20994 18728 20996 18737
rect 21048 18728 21050 18737
rect 20904 18692 20956 18698
rect 20994 18663 21050 18672
rect 20904 18634 20956 18640
rect 20812 18624 20864 18630
rect 20916 18601 20944 18634
rect 20812 18566 20864 18572
rect 20902 18592 20958 18601
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20824 17814 20852 18566
rect 20902 18527 20958 18536
rect 20902 18320 20958 18329
rect 20902 18255 20904 18264
rect 20956 18255 20958 18264
rect 20904 18226 20956 18232
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20720 17672 20772 17678
rect 20772 17632 20852 17660
rect 20720 17614 20772 17620
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20548 16794 20576 16934
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20456 16646 20576 16674
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20352 14952 20404 14958
rect 20272 14912 20352 14940
rect 20352 14894 20404 14900
rect 20364 14074 20392 14894
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20364 13841 20392 13874
rect 20350 13832 20406 13841
rect 20076 13796 20128 13802
rect 20350 13767 20406 13776
rect 20076 13738 20128 13744
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19522 13424 19578 13433
rect 19432 13388 19484 13394
rect 20088 13376 20116 13738
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 19522 13359 19578 13368
rect 19432 13330 19484 13336
rect 19996 13348 20116 13376
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19352 12714 19380 13262
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19246 10704 19302 10713
rect 19246 10639 19248 10648
rect 19300 10639 19302 10648
rect 19248 10610 19300 10616
rect 19352 10554 19380 11494
rect 19260 10526 19380 10554
rect 19444 10554 19472 12786
rect 19996 12170 20024 13348
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 12986 20116 13194
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20272 12850 20300 13670
rect 20350 13424 20406 13433
rect 20350 13359 20406 13368
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20180 11234 20208 12650
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20272 11898 20300 12106
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20180 11206 20300 11234
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19984 10600 20036 10606
rect 19444 10526 19748 10554
rect 19984 10542 20036 10548
rect 19260 9058 19288 10526
rect 19340 10464 19392 10470
rect 19524 10464 19576 10470
rect 19392 10424 19472 10452
rect 19340 10406 19392 10412
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19352 9926 19380 10066
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19352 9178 19380 9522
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19260 9030 19380 9058
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8498 19288 8910
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 7868 19288 8434
rect 19352 7970 19380 9030
rect 19444 8974 19472 10424
rect 19524 10406 19576 10412
rect 19536 10198 19564 10406
rect 19720 10266 19748 10526
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19996 10198 20024 10542
rect 19524 10192 19576 10198
rect 19524 10134 19576 10140
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19536 9217 19564 9590
rect 19996 9353 20024 10134
rect 20088 10130 20116 10610
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20088 9976 20116 10066
rect 20079 9948 20116 9976
rect 20079 9674 20107 9948
rect 20079 9646 20116 9674
rect 19982 9344 20038 9353
rect 19982 9279 20038 9288
rect 19522 9208 19578 9217
rect 19522 9143 19578 9152
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19812 9042 19840 9114
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19996 8974 20024 9279
rect 20088 9178 20116 9646
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19430 8664 19486 8673
rect 19574 8656 19882 8676
rect 19430 8599 19432 8608
rect 19484 8599 19486 8608
rect 19432 8570 19484 8576
rect 19982 8528 20038 8537
rect 19892 8492 19944 8498
rect 19982 8463 20038 8472
rect 19892 8434 19944 8440
rect 19352 7942 19472 7970
rect 19340 7880 19392 7886
rect 19260 7840 19340 7868
rect 19340 7822 19392 7828
rect 19444 7528 19472 7942
rect 19904 7886 19932 8434
rect 19996 8362 20024 8463
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19444 7500 19564 7528
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 5710 19380 7142
rect 19444 7002 19472 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6644 19564 7500
rect 19892 7268 19944 7274
rect 19996 7256 20024 8298
rect 20180 8090 20208 10474
rect 20272 10169 20300 11206
rect 20258 10160 20314 10169
rect 20258 10095 20314 10104
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20272 8838 20300 9862
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20258 8664 20314 8673
rect 20258 8599 20314 8608
rect 20272 8566 20300 8599
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20364 8294 20392 13359
rect 20456 10810 20484 16526
rect 20548 14793 20576 16646
rect 20534 14784 20590 14793
rect 20534 14719 20590 14728
rect 20640 14414 20668 16934
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 15434 20760 16594
rect 20824 15910 20852 17632
rect 20916 17490 20944 18090
rect 21008 17678 21036 18663
rect 21100 18329 21128 18770
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 21192 17882 21220 19479
rect 21284 18426 21312 19654
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21088 17536 21140 17542
rect 20916 17462 21036 17490
rect 21088 17478 21140 17484
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20824 14958 20852 15846
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20824 14226 20852 14894
rect 20916 14346 20944 16934
rect 21008 16522 21036 17462
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 21008 15978 21036 16458
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21008 15473 21036 15506
rect 20994 15464 21050 15473
rect 20994 15399 21050 15408
rect 21100 14929 21128 17478
rect 21086 14920 21142 14929
rect 21086 14855 21142 14864
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21086 14784 21142 14793
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20824 14198 20944 14226
rect 20628 14068 20680 14074
rect 20812 14068 20864 14074
rect 20628 14010 20680 14016
rect 20732 14028 20812 14056
rect 20534 13968 20590 13977
rect 20534 13903 20590 13912
rect 20548 13870 20576 13903
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20548 12730 20576 13806
rect 20640 13190 20668 14010
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20640 12850 20668 13126
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20548 12702 20668 12730
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20456 9586 20484 9930
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20456 9042 20484 9522
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20442 8392 20498 8401
rect 20442 8327 20498 8336
rect 20456 8294 20484 8327
rect 20272 8266 20392 8294
rect 20444 8288 20496 8294
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20272 7936 20300 8266
rect 20444 8230 20496 8236
rect 20180 7908 20300 7936
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19944 7228 20024 7256
rect 19892 7210 19944 7216
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19444 6616 19564 6644
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19444 5370 19472 6616
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19996 6458 20024 6734
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19890 6352 19946 6361
rect 19890 6287 19892 6296
rect 19944 6287 19946 6296
rect 19984 6316 20036 6322
rect 19892 6258 19944 6264
rect 19984 6258 20036 6264
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19154 4040 19210 4049
rect 19154 3975 19210 3984
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18800 2514 18828 2586
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 18892 2446 18920 2790
rect 19168 2774 19196 3975
rect 19260 3058 19288 4082
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19352 3641 19380 3674
rect 19338 3632 19394 3641
rect 19338 3567 19394 3576
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19352 2854 19380 3567
rect 19444 3505 19472 4966
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19616 4208 19668 4214
rect 19614 4176 19616 4185
rect 19668 4176 19670 4185
rect 19614 4111 19670 4120
rect 19708 4072 19760 4078
rect 19996 4026 20024 6258
rect 19708 4014 19760 4020
rect 19522 3904 19578 3913
rect 19522 3839 19578 3848
rect 19430 3496 19486 3505
rect 19536 3466 19564 3839
rect 19720 3738 19748 4014
rect 19904 3998 20024 4026
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 3777 19840 3878
rect 19798 3768 19854 3777
rect 19708 3732 19760 3738
rect 19798 3703 19854 3712
rect 19708 3674 19760 3680
rect 19904 3534 19932 3998
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19430 3431 19486 3440
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19432 3188 19484 3194
rect 19426 3136 19432 3176
rect 19426 3130 19484 3136
rect 19426 3074 19454 3130
rect 19426 3046 19564 3074
rect 19430 2952 19486 2961
rect 19536 2938 19564 3046
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19536 2910 19656 2938
rect 19430 2887 19486 2896
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19076 2746 19196 2774
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 19076 800 19104 2746
rect 19352 2582 19380 2790
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19444 800 19472 2887
rect 19628 2854 19656 2910
rect 19616 2848 19668 2854
rect 19812 2825 19840 2994
rect 19616 2790 19668 2796
rect 19798 2816 19854 2825
rect 19798 2751 19854 2760
rect 20088 2650 20116 7822
rect 20180 4146 20208 7908
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20180 3942 20208 4082
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20272 3890 20300 7754
rect 20442 7440 20498 7449
rect 20548 7410 20576 12582
rect 20640 12374 20668 12702
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20640 11801 20668 12310
rect 20732 12186 20760 14028
rect 20812 14010 20864 14016
rect 20732 12158 20852 12186
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20626 11792 20682 11801
rect 20732 11762 20760 11834
rect 20626 11727 20682 11736
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20626 11520 20682 11529
rect 20626 11455 20682 11464
rect 20640 11286 20668 11455
rect 20824 11354 20852 12158
rect 20916 11354 20944 14198
rect 21008 13841 21036 14758
rect 21086 14719 21142 14728
rect 20994 13832 21050 13841
rect 20994 13767 21050 13776
rect 20994 13560 21050 13569
rect 20994 13495 20996 13504
rect 21048 13495 21050 13504
rect 20996 13466 21048 13472
rect 21008 12782 21036 13466
rect 21100 12986 21128 14719
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20996 12776 21048 12782
rect 21048 12736 21128 12764
rect 20996 12718 21048 12724
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20628 11280 20680 11286
rect 21008 11234 21036 11766
rect 20628 11222 20680 11228
rect 20640 8430 20668 11222
rect 20824 11206 21036 11234
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20732 9994 20760 10542
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20732 8378 20760 9930
rect 20824 9330 20852 11206
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20916 9450 20944 10610
rect 21008 10538 21036 11086
rect 21100 11082 21128 12736
rect 21192 12714 21220 17546
rect 21284 17270 21312 18158
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21376 16454 21404 20046
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21456 19848 21508 19854
rect 21454 19816 21456 19825
rect 21508 19816 21510 19825
rect 21454 19751 21510 19760
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 16776 21496 19654
rect 21560 19378 21588 24210
rect 21836 23882 21864 24346
rect 22020 24206 22048 24704
rect 22204 24274 22232 26522
rect 22388 24732 22416 27338
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22572 26994 22600 27270
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22572 26382 22600 26930
rect 24228 26926 24256 27814
rect 24412 27606 24440 28018
rect 24768 27872 24820 27878
rect 24820 27832 24900 27860
rect 24768 27814 24820 27820
rect 24400 27600 24452 27606
rect 24400 27542 24452 27548
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 24216 26920 24268 26926
rect 24216 26862 24268 26868
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 22652 26512 22704 26518
rect 22652 26454 22704 26460
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22572 25906 22600 26318
rect 22664 26246 22692 26454
rect 23112 26308 23164 26314
rect 23112 26250 23164 26256
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 22652 26240 22704 26246
rect 22652 26182 22704 26188
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22664 25786 22692 26182
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22572 25758 22692 25786
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 25362 22508 25638
rect 22572 25362 22600 25758
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 22480 24750 22508 25298
rect 22296 24704 22416 24732
rect 22468 24744 22520 24750
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 21836 23866 21956 23882
rect 21836 23860 21968 23866
rect 21836 23854 21916 23860
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21744 22930 21772 23666
rect 21836 23526 21864 23854
rect 21916 23802 21968 23808
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21824 23112 21876 23118
rect 21928 23066 21956 23598
rect 21876 23060 21956 23066
rect 21824 23054 21956 23060
rect 21836 23038 21956 23054
rect 21744 22902 21864 22930
rect 21836 22642 21864 22902
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21836 21622 21864 22578
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 21638 20632 21694 20641
rect 21638 20567 21640 20576
rect 21692 20567 21694 20576
rect 21640 20538 21692 20544
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21652 18873 21680 20402
rect 21638 18864 21694 18873
rect 21548 18828 21600 18834
rect 21638 18799 21694 18808
rect 21548 18770 21600 18776
rect 21560 17066 21588 18770
rect 21652 18766 21680 18799
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21640 17604 21692 17610
rect 21744 17592 21772 20402
rect 21836 19718 21864 21082
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21836 18601 21864 19382
rect 21822 18592 21878 18601
rect 21822 18527 21878 18536
rect 21928 18408 21956 23038
rect 22020 21622 22048 24142
rect 22204 23730 22232 24210
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21692 17564 21772 17592
rect 21836 18380 21956 18408
rect 21640 17546 21692 17552
rect 21548 17060 21600 17066
rect 21548 17002 21600 17008
rect 21468 16748 21588 16776
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21362 16280 21418 16289
rect 21362 16215 21418 16224
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 13326 21312 14962
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21192 11830 21220 12038
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21086 10976 21142 10985
rect 21086 10911 21142 10920
rect 21100 10674 21128 10911
rect 21192 10674 21220 11222
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21008 10062 21036 10474
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21100 9994 21128 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 21192 9654 21220 9998
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21100 9518 21128 9590
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20824 9302 21128 9330
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 21008 8974 21036 9114
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20824 8673 20852 8842
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20994 8800 21050 8809
rect 20810 8664 20866 8673
rect 20810 8599 20866 8608
rect 20916 8498 20944 8774
rect 20994 8735 21050 8744
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20732 8350 20852 8378
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20442 7375 20498 7384
rect 20536 7404 20588 7410
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20364 6322 20392 6598
rect 20456 6458 20484 7375
rect 20536 7346 20588 7352
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20548 6458 20576 6666
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20364 5914 20392 6258
rect 20534 6216 20590 6225
rect 20444 6180 20496 6186
rect 20534 6151 20590 6160
rect 20444 6122 20496 6128
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20456 5098 20484 6122
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20364 4049 20392 4490
rect 20456 4282 20484 4558
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20350 4040 20406 4049
rect 20350 3975 20406 3984
rect 20272 3862 20484 3890
rect 20258 3632 20314 3641
rect 20258 3567 20314 3576
rect 20352 3596 20404 3602
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19522 2544 19578 2553
rect 19522 2479 19578 2488
rect 19536 2446 19564 2479
rect 20180 2446 20208 3334
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19812 800 19840 1906
rect 20272 1170 20300 3567
rect 20352 3538 20404 3544
rect 20364 3126 20392 3538
rect 20456 3210 20484 3862
rect 20548 3534 20576 6151
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20456 3182 20576 3210
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20548 3058 20576 3182
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20456 1902 20484 2994
rect 20534 2952 20590 2961
rect 20534 2887 20590 2896
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20180 1142 20300 1170
rect 20180 800 20208 1142
rect 20548 800 20576 2887
rect 20640 2650 20668 7822
rect 20732 7698 20760 8230
rect 20824 7818 20852 8350
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20732 7670 20852 7698
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20732 5234 20760 6666
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20824 5166 20852 7670
rect 21008 6866 21036 8735
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20994 6624 21050 6633
rect 20994 6559 21050 6568
rect 21008 6361 21036 6559
rect 20994 6352 21050 6361
rect 20994 6287 20996 6296
rect 21048 6287 21050 6296
rect 20996 6258 21048 6264
rect 21008 6227 21036 6258
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 20718 4176 20774 4185
rect 20718 4111 20720 4120
rect 20772 4111 20774 4120
rect 20720 4082 20772 4088
rect 20732 3534 20760 4082
rect 20824 3641 20852 4422
rect 20810 3632 20866 3641
rect 20810 3567 20866 3576
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20824 3194 20852 3402
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20640 1426 20668 2246
rect 20628 1420 20680 1426
rect 20628 1362 20680 1368
rect 20916 800 20944 4422
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 21008 4049 21036 4082
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 21008 2854 21036 3470
rect 21100 2990 21128 9302
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21192 8838 21220 8910
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21284 8294 21312 12786
rect 21376 9178 21404 16215
rect 21468 15502 21496 16594
rect 21560 16590 21588 16748
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 16425 21588 16526
rect 21546 16416 21602 16425
rect 21546 16351 21602 16360
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21560 16017 21588 16186
rect 21652 16114 21680 17546
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21744 16969 21772 17070
rect 21730 16960 21786 16969
rect 21730 16895 21786 16904
rect 21730 16824 21786 16833
rect 21730 16759 21786 16768
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21546 16008 21602 16017
rect 21546 15943 21602 15952
rect 21546 15600 21602 15609
rect 21546 15535 21602 15544
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 14890 21496 15438
rect 21560 15162 21588 15535
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21468 12434 21496 14826
rect 21546 14648 21602 14657
rect 21546 14583 21602 14592
rect 21560 14414 21588 14583
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21744 13938 21772 16759
rect 21836 15638 21864 18380
rect 22020 18290 22048 21558
rect 22112 19990 22140 22646
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 19990 22232 20742
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22112 18970 22140 19790
rect 22204 19514 22232 19790
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18306 22232 18566
rect 22296 18426 22324 24704
rect 22468 24686 22520 24692
rect 22572 24562 22600 25298
rect 22480 24534 22600 24562
rect 22480 24274 22508 24534
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22388 22710 22416 22918
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22480 22094 22508 24210
rect 22756 23712 22784 25910
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22848 24682 22876 25842
rect 23124 25838 23152 26250
rect 23112 25832 23164 25838
rect 23112 25774 23164 25780
rect 23020 25356 23072 25362
rect 23020 25298 23072 25304
rect 23032 24818 23060 25298
rect 23124 25294 23152 25774
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 24313 23520 24550
rect 23478 24304 23534 24313
rect 23478 24239 23534 24248
rect 22836 23724 22888 23730
rect 22756 23684 22836 23712
rect 22836 23666 22888 23672
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 22438 22600 23462
rect 22926 23352 22982 23361
rect 22926 23287 22928 23296
rect 22980 23287 22982 23296
rect 22928 23258 22980 23264
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22388 22066 22508 22094
rect 22388 20448 22416 22066
rect 22572 21554 22600 22374
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 23032 21622 23060 21898
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22650 21448 22706 21457
rect 22650 21383 22706 21392
rect 22664 21078 22692 21383
rect 22652 21072 22704 21078
rect 22652 21014 22704 21020
rect 22744 21072 22796 21078
rect 22744 21014 22796 21020
rect 22664 20602 22692 21014
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22388 20420 22692 20448
rect 22374 19952 22430 19961
rect 22374 19887 22430 19896
rect 22388 19854 22416 19887
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22468 18760 22520 18766
rect 22466 18728 22468 18737
rect 22520 18728 22522 18737
rect 22466 18663 22522 18672
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22008 18284 22060 18290
rect 22204 18278 22324 18306
rect 22008 18226 22060 18232
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16017 21956 16934
rect 21914 16008 21970 16017
rect 22098 16008 22154 16017
rect 21914 15943 21970 15952
rect 22008 15972 22060 15978
rect 22098 15943 22154 15952
rect 22008 15914 22060 15920
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15026 21864 15438
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21836 13818 21864 14962
rect 21744 13790 21864 13818
rect 21744 13297 21772 13790
rect 21730 13288 21786 13297
rect 21730 13223 21786 13232
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21468 12406 21588 12434
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 11150 21496 11630
rect 21560 11286 21588 12406
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21468 10606 21496 11086
rect 21560 10674 21588 11086
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21468 10130 21496 10542
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21454 10024 21510 10033
rect 21454 9959 21510 9968
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21376 8090 21404 8230
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 3466 21220 7686
rect 21284 7546 21312 7822
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 4758 21312 6258
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21284 1970 21312 4150
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 21376 1834 21404 4966
rect 21468 3398 21496 9959
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21468 1970 21496 2994
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 21364 1828 21416 1834
rect 21364 1770 21416 1776
rect 21284 870 21404 898
rect 21284 800 21312 870
rect 14752 734 14964 762
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21376 762 21404 870
rect 21560 762 21588 10202
rect 21652 7818 21680 12718
rect 21744 11218 21772 13223
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21730 10976 21786 10985
rect 21730 10911 21786 10920
rect 21744 9586 21772 10911
rect 21836 9625 21864 11018
rect 21928 10742 21956 15846
rect 22020 15162 22048 15914
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22112 15094 22140 15943
rect 22204 15910 22232 17206
rect 22296 17134 22324 18278
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22190 14648 22246 14657
rect 22296 14618 22324 17070
rect 22190 14583 22246 14592
rect 22284 14612 22336 14618
rect 22098 14512 22154 14521
rect 22098 14447 22154 14456
rect 22112 14414 22140 14447
rect 22204 14414 22232 14583
rect 22284 14554 22336 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22008 14272 22060 14278
rect 22006 14240 22008 14249
rect 22060 14240 22062 14249
rect 22006 14175 22062 14184
rect 22008 13932 22060 13938
rect 22112 13920 22140 14350
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 14006 22232 14214
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22060 13892 22140 13920
rect 22008 13874 22060 13880
rect 22020 12850 22048 13874
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22020 11762 22048 12786
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22020 10674 22048 11562
rect 22112 11082 22140 13330
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12753 22232 13262
rect 22190 12744 22246 12753
rect 22190 12679 22246 12688
rect 22296 12356 22324 14554
rect 22388 12458 22416 18022
rect 22480 17746 22508 18362
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22572 17116 22600 19246
rect 22664 18222 22692 20420
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22664 17270 22692 17478
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22652 17128 22704 17134
rect 22572 17088 22652 17116
rect 22652 17070 22704 17076
rect 22664 16114 22692 17070
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22756 15892 22784 21014
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 19378 22876 20742
rect 23124 20466 23152 21966
rect 23216 21486 23244 23054
rect 23584 22982 23612 26250
rect 23768 25294 23796 26726
rect 23860 26586 23888 26862
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 24044 26586 24072 26794
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 24228 26518 24256 26862
rect 24216 26512 24268 26518
rect 24216 26454 24268 26460
rect 24308 25900 24360 25906
rect 24308 25842 24360 25848
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23768 23186 23796 24890
rect 23848 23588 23900 23594
rect 23848 23530 23900 23536
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23756 23044 23808 23050
rect 23756 22986 23808 22992
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23768 22438 23796 22986
rect 23860 22982 23888 23530
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23860 22506 23888 22918
rect 23848 22500 23900 22506
rect 23848 22442 23900 22448
rect 23756 22432 23808 22438
rect 23808 22380 23888 22386
rect 23756 22374 23888 22380
rect 23768 22358 23888 22374
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21554 23520 21830
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23216 21078 23244 21422
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22836 19372 22888 19378
rect 23124 19334 23152 20198
rect 22836 19314 22888 19320
rect 23032 19306 23152 19334
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22940 18290 22968 18634
rect 23032 18426 23060 19306
rect 23216 18698 23244 20538
rect 23308 18970 23336 21014
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23400 20058 23428 20402
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23492 19854 23520 20878
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23204 18692 23256 18698
rect 23256 18652 23336 18680
rect 23204 18634 23256 18640
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22572 15864 22784 15892
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 14550 22508 15302
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22480 14385 22508 14486
rect 22466 14376 22522 14385
rect 22466 14311 22522 14320
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22480 13326 22508 13738
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12986 22508 13126
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22480 12617 22508 12718
rect 22466 12608 22522 12617
rect 22466 12543 22522 12552
rect 22388 12430 22508 12458
rect 22296 12328 22416 12356
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22112 10538 22140 11018
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 21916 9716 21968 9722
rect 22204 9674 22232 11494
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 21916 9658 21968 9664
rect 21822 9616 21878 9625
rect 21732 9580 21784 9586
rect 21822 9551 21878 9560
rect 21732 9522 21784 9528
rect 21744 8906 21772 9522
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21836 8945 21864 9046
rect 21822 8936 21878 8945
rect 21732 8900 21784 8906
rect 21928 8906 21956 9658
rect 22020 9646 22232 9674
rect 22296 9654 22324 11154
rect 22388 9722 22416 12328
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 9648 22336 9654
rect 22020 9081 22048 9646
rect 22284 9590 22336 9596
rect 22374 9616 22430 9625
rect 22374 9551 22430 9560
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22100 9376 22152 9382
rect 22098 9344 22100 9353
rect 22192 9376 22244 9382
rect 22152 9344 22154 9353
rect 22192 9318 22244 9324
rect 22098 9279 22154 9288
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 22204 8974 22232 9318
rect 22296 9178 22324 9454
rect 22388 9178 22416 9551
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 21822 8871 21878 8880
rect 21916 8900 21968 8906
rect 21732 8842 21784 8848
rect 21916 8842 21968 8848
rect 21744 8566 21772 8842
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21836 8634 21864 8774
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21744 5574 21772 8502
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22020 8401 22048 8434
rect 22006 8392 22062 8401
rect 22006 8327 22062 8336
rect 22480 8294 22508 12430
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 22204 8266 22508 8294
rect 21836 7954 21864 8230
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 22020 7410 22048 7754
rect 22112 7478 22140 7822
rect 22100 7472 22152 7478
rect 22100 7414 22152 7420
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22020 5710 22048 6734
rect 22112 6322 22140 6802
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21652 800 21680 2790
rect 22204 2530 22232 8266
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22296 6798 22324 7210
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22388 6361 22416 7414
rect 22572 6746 22600 15864
rect 22650 15736 22706 15745
rect 22650 15671 22706 15680
rect 22664 14958 22692 15671
rect 22848 15638 22876 18158
rect 23032 18086 23060 18158
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 23124 17898 23152 18566
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23032 17870 23152 17898
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 16998 22968 17614
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14414 22692 14758
rect 22940 14464 22968 16526
rect 22848 14436 22968 14464
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22744 14408 22796 14414
rect 22848 14396 22876 14436
rect 22796 14368 22876 14396
rect 22744 14350 22796 14356
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22664 9625 22692 13806
rect 22756 12764 22784 13806
rect 22848 12918 22876 13874
rect 22940 13870 22968 14282
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 23032 13802 23060 17870
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 23124 17678 23152 17750
rect 23216 17746 23244 18158
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23216 17270 23244 17682
rect 23308 17678 23336 18652
rect 23388 18080 23440 18086
rect 23386 18048 23388 18057
rect 23440 18048 23442 18057
rect 23386 17983 23442 17992
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23216 16590 23244 17206
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23216 16046 23244 16526
rect 23308 16250 23336 16526
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23110 14512 23166 14521
rect 23110 14447 23166 14456
rect 23124 14414 23152 14447
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23124 13530 23152 14350
rect 23216 13802 23244 14758
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22756 12736 22876 12764
rect 22742 12608 22798 12617
rect 22742 12543 22798 12552
rect 22756 12238 22784 12543
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22848 11898 22876 12736
rect 22940 12730 22968 13330
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12850 23060 13126
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22940 12702 23060 12730
rect 23032 12434 23060 12702
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 22940 12406 23060 12434
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22834 11792 22890 11801
rect 22834 11727 22890 11736
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22664 9081 22692 9114
rect 22650 9072 22706 9081
rect 22650 9007 22706 9016
rect 22664 8362 22692 9007
rect 22756 8906 22784 10474
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22664 7002 22692 8298
rect 22848 7750 22876 11727
rect 22940 10305 22968 12406
rect 23124 12238 23152 12582
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23110 11656 23166 11665
rect 23110 11591 23166 11600
rect 23124 11150 23152 11591
rect 23216 11354 23244 12038
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23202 11248 23258 11257
rect 23202 11183 23258 11192
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23216 11014 23244 11183
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 23216 10606 23244 10950
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 22926 10296 22982 10305
rect 22926 10231 22982 10240
rect 22926 10160 22982 10169
rect 22926 10095 22982 10104
rect 22836 7744 22888 7750
rect 22940 7721 22968 10095
rect 23216 9674 23244 10542
rect 23124 9646 23244 9674
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 9178 23060 9318
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 8566 23060 8910
rect 23124 8634 23152 9646
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23020 8424 23072 8430
rect 23018 8392 23020 8401
rect 23072 8392 23074 8401
rect 23018 8327 23074 8336
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 22836 7686 22888 7692
rect 22926 7712 22982 7721
rect 22926 7647 22982 7656
rect 23032 7546 23060 8230
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22480 6718 22600 6746
rect 22652 6792 22704 6798
rect 22704 6752 22784 6780
rect 22652 6734 22704 6740
rect 22480 6458 22508 6718
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22374 6352 22430 6361
rect 22374 6287 22376 6296
rect 22428 6287 22430 6296
rect 22376 6258 22428 6264
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22296 5030 22324 5170
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22296 2854 22324 4422
rect 22388 4146 22416 6258
rect 22572 5370 22600 6598
rect 22756 6458 22784 6752
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22664 5098 22692 6258
rect 22756 5846 22784 6394
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22756 5234 22784 5510
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22480 4978 22508 5034
rect 22480 4950 22600 4978
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22388 3738 22416 4082
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22480 2774 22508 4422
rect 22572 4282 22600 4950
rect 22848 4622 22876 7142
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22940 5710 22968 6666
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 23032 3534 23060 7482
rect 23124 6934 23152 8570
rect 23308 8401 23336 14214
rect 23400 13734 23428 16662
rect 23492 15026 23520 19654
rect 23584 19378 23612 20742
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23584 18902 23612 19314
rect 23676 18902 23704 21354
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23768 21146 23796 21286
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23664 18896 23716 18902
rect 23664 18838 23716 18844
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23584 16590 23612 17614
rect 23676 16794 23704 18838
rect 23768 18766 23796 19110
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23584 15162 23612 15914
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 14249 23520 14758
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23478 14240 23534 14249
rect 23478 14175 23534 14184
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23492 12322 23520 12922
rect 23400 12294 23520 12322
rect 23400 12238 23428 12294
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23400 11150 23428 11698
rect 23492 11354 23520 12106
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23386 10296 23442 10305
rect 23386 10231 23442 10240
rect 23294 8392 23350 8401
rect 23294 8327 23350 8336
rect 23294 7304 23350 7313
rect 23400 7274 23428 10231
rect 23492 10062 23520 11290
rect 23584 10985 23612 14554
rect 23768 12918 23796 18702
rect 23860 14346 23888 22358
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23952 12434 23980 25162
rect 24320 24818 24348 25842
rect 24596 25498 24624 27406
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 24044 24206 24072 24550
rect 24228 24410 24256 24754
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 24030 23488 24086 23497
rect 24030 23423 24086 23432
rect 24044 23186 24072 23423
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24044 19174 24072 23122
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 24044 18834 24072 19110
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24032 16992 24084 16998
rect 24136 16980 24164 24210
rect 24688 24206 24716 26318
rect 24780 25838 24808 26862
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24780 25498 24808 25774
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24872 25362 24900 27832
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24780 23866 24808 24754
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24320 23526 24348 23802
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24228 21570 24256 21898
rect 24320 21690 24348 23462
rect 24780 23186 24808 23462
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24872 23118 24900 25298
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24308 21684 24360 21690
rect 24308 21626 24360 21632
rect 24228 21542 24348 21570
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 24084 16952 24164 16980
rect 24032 16934 24084 16940
rect 24044 13705 24072 16934
rect 24228 15858 24256 20810
rect 24320 20262 24348 21542
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24320 19718 24348 20198
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 24320 16658 24348 17002
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24412 16232 24440 22170
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24492 21956 24544 21962
rect 24492 21898 24544 21904
rect 24504 19990 24532 21898
rect 24596 20058 24624 22034
rect 24872 22030 24900 23054
rect 24964 22930 24992 35866
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 25056 26466 25084 26726
rect 25148 26586 25176 28018
rect 26056 27872 26108 27878
rect 26056 27814 26108 27820
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25240 27062 25268 27406
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25240 26858 25268 26998
rect 25228 26852 25280 26858
rect 25228 26794 25280 26800
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25228 26512 25280 26518
rect 25056 26438 25176 26466
rect 25228 26454 25280 26460
rect 25148 25294 25176 26438
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 25056 23662 25084 25162
rect 25148 24954 25176 25230
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25240 24682 25268 26454
rect 25332 26382 25360 27270
rect 26068 26994 26096 27814
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 26240 27056 26292 27062
rect 26240 26998 26292 27004
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25608 26382 25636 26726
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25332 25906 25360 25978
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25412 25764 25464 25770
rect 25412 25706 25464 25712
rect 25228 24676 25280 24682
rect 25228 24618 25280 24624
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25044 23656 25096 23662
rect 25096 23616 25176 23644
rect 25044 23598 25096 23604
rect 24964 22902 25084 22930
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24492 19984 24544 19990
rect 24492 19926 24544 19932
rect 24504 19446 24532 19926
rect 24688 19786 24716 20334
rect 24780 19802 24808 21354
rect 24872 21010 24900 21490
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24872 20466 24900 20946
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24860 19848 24912 19854
rect 24780 19796 24860 19802
rect 24780 19790 24912 19796
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24780 19774 24900 19790
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24584 18692 24636 18698
rect 24584 18634 24636 18640
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24504 17202 24532 18226
rect 24596 18154 24624 18634
rect 24688 18290 24716 19722
rect 24780 19378 24808 19774
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24964 19281 24992 22578
rect 25056 19514 25084 22902
rect 25148 21146 25176 23616
rect 25228 23588 25280 23594
rect 25228 23530 25280 23536
rect 25240 23497 25268 23530
rect 25226 23488 25282 23497
rect 25226 23423 25282 23432
rect 25332 22137 25360 23734
rect 25318 22128 25374 22137
rect 25318 22063 25374 22072
rect 25332 21350 25360 22063
rect 25424 21690 25452 25706
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25700 25294 25728 25638
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25608 24070 25636 24686
rect 25792 24154 25820 26318
rect 25700 24126 25820 24154
rect 26068 24138 26096 26930
rect 26252 26382 26280 26998
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26424 26852 26476 26858
rect 26424 26794 26476 26800
rect 26436 26382 26464 26794
rect 26896 26586 26924 26930
rect 27620 26784 27672 26790
rect 27620 26726 27672 26732
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 26240 26376 26292 26382
rect 26424 26376 26476 26382
rect 26292 26336 26372 26364
rect 26240 26318 26292 26324
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26252 25158 26280 25842
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 24954 26280 25094
rect 26240 24948 26292 24954
rect 26240 24890 26292 24896
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 26056 24132 26108 24138
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25700 23798 25728 24126
rect 26056 24074 26108 24080
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25688 23792 25740 23798
rect 25688 23734 25740 23740
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25516 23361 25544 23666
rect 25502 23352 25558 23361
rect 25502 23287 25558 23296
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25516 22098 25544 22510
rect 25608 22234 25636 23054
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25136 21140 25188 21146
rect 25188 21100 25268 21128
rect 25136 21082 25188 21088
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24950 19272 25006 19281
rect 24950 19207 25006 19216
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24596 17338 24624 17546
rect 24688 17338 24716 18226
rect 24872 18154 24900 18566
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24964 17678 24992 18022
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24780 17202 24808 17478
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24872 16794 24900 17614
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25056 16969 25084 17138
rect 25042 16960 25098 16969
rect 25042 16895 25098 16904
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24674 16552 24730 16561
rect 24674 16487 24730 16496
rect 24412 16204 24532 16232
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24228 15830 24348 15858
rect 24320 15144 24348 15830
rect 24412 15706 24440 16050
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24320 15116 24440 15144
rect 24214 15056 24270 15065
rect 24214 14991 24216 15000
rect 24268 14991 24270 15000
rect 24216 14962 24268 14968
rect 24124 14952 24176 14958
rect 24122 14920 24124 14929
rect 24176 14920 24178 14929
rect 24122 14855 24178 14864
rect 24030 13696 24086 13705
rect 24030 13631 24086 13640
rect 24228 13462 24256 14962
rect 24412 14822 24440 15116
rect 24504 15008 24532 16204
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24596 15366 24624 15506
rect 24688 15502 24716 16487
rect 24872 16182 24900 16730
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24872 15620 24900 16118
rect 24964 15881 24992 16118
rect 24950 15872 25006 15881
rect 24950 15807 25006 15816
rect 25044 15632 25096 15638
rect 24872 15592 25044 15620
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24676 15020 24728 15026
rect 24504 14980 24676 15008
rect 24400 14816 24452 14822
rect 24398 14784 24400 14793
rect 24452 14784 24454 14793
rect 24398 14719 24454 14728
rect 24412 14693 24440 14719
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24136 12753 24164 13330
rect 24122 12744 24178 12753
rect 24122 12679 24124 12688
rect 24176 12679 24178 12688
rect 24124 12650 24176 12656
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 23768 12406 23980 12434
rect 23570 10976 23626 10985
rect 23570 10911 23626 10920
rect 23768 10826 23796 12406
rect 24228 12374 24256 12582
rect 24216 12368 24268 12374
rect 24216 12310 24268 12316
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 11898 24072 12174
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23860 11150 23888 11766
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23584 10798 23796 10826
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23492 8090 23520 8434
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23294 7239 23350 7248
rect 23388 7268 23440 7274
rect 23308 6934 23336 7239
rect 23388 7210 23440 7216
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 23308 5574 23336 6870
rect 23584 6798 23612 10798
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23938 10704 23994 10713
rect 23676 10538 23704 10678
rect 23756 10668 23808 10674
rect 23938 10639 23994 10648
rect 23756 10610 23808 10616
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23768 10266 23796 10610
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23860 10146 23888 10406
rect 23768 10118 23888 10146
rect 23768 9654 23796 10118
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23676 8974 23704 9454
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23478 6080 23534 6089
rect 23478 6015 23534 6024
rect 23386 5944 23442 5953
rect 23492 5914 23520 6015
rect 23386 5879 23388 5888
rect 23440 5879 23442 5888
rect 23480 5908 23532 5914
rect 23388 5850 23440 5856
rect 23480 5850 23532 5856
rect 23584 5778 23612 6190
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23388 5704 23440 5710
rect 23676 5658 23704 7890
rect 23388 5646 23440 5652
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23308 5234 23336 5510
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23308 3913 23336 3946
rect 23400 3924 23428 5646
rect 23584 5630 23704 5658
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4146 23520 4966
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23480 3936 23532 3942
rect 23294 3904 23350 3913
rect 23400 3896 23480 3924
rect 23480 3878 23532 3884
rect 23294 3839 23350 3848
rect 23492 3777 23520 3878
rect 23478 3768 23534 3777
rect 23478 3703 23534 3712
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22112 2502 22232 2530
rect 22388 2746 22508 2774
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22020 800 22048 2382
rect 22112 1766 22140 2502
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22204 2106 22232 2382
rect 22192 2100 22244 2106
rect 22192 2042 22244 2048
rect 22100 1760 22152 1766
rect 22100 1702 22152 1708
rect 22388 800 22416 2746
rect 22756 800 22784 2858
rect 23124 800 23152 3606
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23308 2514 23336 3334
rect 23400 3058 23428 3538
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23492 2990 23520 3402
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23584 2774 23612 5630
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23676 5234 23704 5510
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23768 5114 23796 9590
rect 23860 6882 23888 9930
rect 23952 7954 23980 10639
rect 24030 9616 24086 9625
rect 24030 9551 24086 9560
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 24044 7410 24072 9551
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24136 8022 24164 8434
rect 24228 8362 24256 12310
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24228 7886 24256 8298
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23952 7290 23980 7346
rect 24320 7324 24348 14010
rect 24412 13326 24440 14350
rect 24504 13530 24532 14980
rect 24676 14962 24728 14968
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24596 14074 24624 14758
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24688 13802 24716 14350
rect 24780 14346 24808 15574
rect 24872 15026 24900 15592
rect 25044 15574 25096 15580
rect 24950 15192 25006 15201
rect 24950 15127 25006 15136
rect 24964 15094 24992 15127
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24858 14784 24914 14793
rect 24858 14719 24914 14728
rect 24872 14362 24900 14719
rect 25056 14414 25084 14826
rect 25044 14408 25096 14414
rect 24768 14340 24820 14346
rect 24872 14334 24992 14362
rect 25044 14350 25096 14356
rect 24768 14282 24820 14288
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 13938 24900 14214
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24676 13796 24728 13802
rect 24676 13738 24728 13744
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24688 13326 24716 13738
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24412 12850 24440 13262
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 8838 24440 12786
rect 24688 12714 24716 13262
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24504 11830 24532 12174
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24584 11620 24636 11626
rect 24504 11580 24584 11608
rect 24504 10606 24532 11580
rect 24584 11562 24636 11568
rect 24688 11218 24716 12650
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24504 9042 24532 9998
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24596 8090 24624 11018
rect 24674 9616 24730 9625
rect 24674 9551 24676 9560
rect 24728 9551 24730 9560
rect 24676 9522 24728 9528
rect 24688 8566 24716 9522
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24596 7478 24624 8026
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24688 7546 24716 7754
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24780 7410 24808 13398
rect 24872 13326 24900 13738
rect 24964 13394 24992 14334
rect 25148 13802 25176 19926
rect 25240 18902 25268 21100
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25332 20210 25360 20878
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 25516 20398 25544 20810
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25608 20330 25636 21558
rect 25700 21554 25728 22442
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25332 20182 25544 20210
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25240 18358 25268 18838
rect 25332 18834 25360 19654
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25320 18828 25372 18834
rect 25320 18770 25372 18776
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25332 18290 25360 18566
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 17218 25360 18226
rect 25424 17338 25452 19314
rect 25516 18154 25544 20182
rect 25700 19700 25728 21490
rect 25792 21146 25820 24006
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25884 22030 25912 22646
rect 25976 22438 26004 23666
rect 26160 23322 26188 24822
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26252 24410 26280 24754
rect 26344 24682 26372 26336
rect 26424 26318 26476 26324
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26516 26308 26568 26314
rect 26516 26250 26568 26256
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26528 24614 26556 26250
rect 27080 26042 27108 26318
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26804 24818 26832 25774
rect 27172 25226 27200 25842
rect 27632 25294 27660 26726
rect 27908 26382 27936 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27988 26376 28040 26382
rect 27988 26318 28040 26324
rect 27724 25838 27752 26318
rect 27804 26308 27856 26314
rect 27804 26250 27856 26256
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27160 25220 27212 25226
rect 27160 25162 27212 25168
rect 27632 24954 27660 25230
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 26068 22574 26096 22918
rect 26160 22642 26188 23258
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26056 22568 26108 22574
rect 26056 22510 26108 22516
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 25976 22234 26004 22374
rect 25964 22228 26016 22234
rect 25964 22170 26016 22176
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25884 21434 25912 21966
rect 25976 21622 26004 22170
rect 26160 22094 26188 22578
rect 26988 22166 27016 24754
rect 27632 24732 27660 24890
rect 27724 24818 27752 25774
rect 27816 25770 27844 26250
rect 28000 25922 28028 26318
rect 28080 26240 28132 26246
rect 28080 26182 28132 26188
rect 27908 25906 28028 25922
rect 28092 25906 28120 26182
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 27896 25900 28028 25906
rect 27948 25894 28028 25900
rect 28080 25900 28132 25906
rect 27896 25842 27948 25848
rect 28080 25842 28132 25848
rect 28264 25900 28316 25906
rect 28264 25842 28316 25848
rect 27804 25764 27856 25770
rect 27804 25706 27856 25712
rect 27896 25696 27948 25702
rect 27896 25638 27948 25644
rect 27908 25294 27936 25638
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 28172 25152 28224 25158
rect 28172 25094 28224 25100
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27356 24704 27660 24732
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27080 23254 27108 24550
rect 27068 23248 27120 23254
rect 27068 23190 27120 23196
rect 27160 23044 27212 23050
rect 27160 22986 27212 22992
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26160 22066 26280 22094
rect 26252 22030 26280 22066
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26332 21888 26384 21894
rect 26332 21830 26384 21836
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 25964 21480 26016 21486
rect 25884 21428 25964 21434
rect 25884 21422 26016 21428
rect 25884 21406 26004 21422
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25792 19854 25820 21082
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25700 19672 25820 19700
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25504 18148 25556 18154
rect 25504 18090 25556 18096
rect 25608 18034 25636 18362
rect 25516 18006 25636 18034
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25332 17202 25452 17218
rect 25332 17196 25464 17202
rect 25332 17190 25412 17196
rect 25412 17138 25464 17144
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 16250 25268 16526
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25332 15502 25360 17070
rect 25424 15910 25452 17138
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25332 14929 25360 14962
rect 25318 14920 25374 14929
rect 25318 14855 25374 14864
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24872 12102 24900 12650
rect 25056 12442 25084 12650
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24860 11688 24912 11694
rect 25056 11642 25084 12378
rect 24912 11636 25084 11642
rect 24860 11630 25084 11636
rect 24872 11614 25084 11630
rect 25056 11558 25084 11614
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24872 10674 24900 11290
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24872 9518 24900 10610
rect 24964 9586 24992 11494
rect 25148 9674 25176 13738
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25240 12782 25268 13670
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25332 12646 25360 13670
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25240 11830 25268 12038
rect 25424 11898 25452 15846
rect 25516 12918 25544 18006
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25608 16590 25636 17546
rect 25792 16726 25820 19672
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25884 18698 25912 19246
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25884 18290 25912 18634
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25884 17542 25912 18226
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25780 16720 25832 16726
rect 25780 16662 25832 16668
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25608 15502 25636 16390
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25700 15348 25728 16594
rect 25608 15320 25728 15348
rect 25608 15162 25636 15320
rect 25686 15192 25742 15201
rect 25596 15156 25648 15162
rect 25686 15127 25742 15136
rect 25596 15098 25648 15104
rect 25608 14550 25636 15098
rect 25700 15094 25728 15127
rect 25688 15088 25740 15094
rect 25688 15030 25740 15036
rect 25792 14618 25820 16662
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 13870 25728 14214
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25686 13696 25742 13705
rect 25686 13631 25742 13640
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25608 12434 25636 13262
rect 25700 12918 25728 13631
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25608 12406 25728 12434
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25608 11218 25636 12038
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25502 11112 25558 11121
rect 25502 11047 25558 11056
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25240 9722 25268 10542
rect 25139 9646 25176 9674
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25139 9602 25167 9646
rect 24952 9580 25004 9586
rect 25139 9574 25176 9602
rect 24952 9522 25004 9528
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 25042 8664 25098 8673
rect 25042 8599 25044 8608
rect 25096 8599 25098 8608
rect 25044 8570 25096 8576
rect 24952 8356 25004 8362
rect 24872 8316 24952 8344
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24320 7296 24624 7324
rect 23952 7262 24164 7290
rect 23860 6854 23980 6882
rect 23676 5086 23796 5114
rect 23676 3058 23704 5086
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 3670 23796 4422
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23492 2746 23612 2774
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23492 800 23520 2746
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23860 800 23888 2246
rect 21376 734 21588 762
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 23952 762 23980 6854
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24044 6118 24072 6394
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4214 24072 5102
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 24136 3398 24164 7262
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24320 6798 24348 7142
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24320 6361 24348 6734
rect 24306 6352 24362 6361
rect 24306 6287 24362 6296
rect 24320 5710 24348 6287
rect 24412 6186 24440 7142
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 3534 24256 4422
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24044 3126 24072 3334
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 24228 2990 24256 3470
rect 24320 3194 24348 5170
rect 24412 4146 24440 6122
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24504 5642 24532 6054
rect 24492 5636 24544 5642
rect 24492 5578 24544 5584
rect 24596 5522 24624 7296
rect 24872 6610 24900 8316
rect 24952 8298 25004 8304
rect 25148 8022 25176 9574
rect 25417 9564 25469 9570
rect 25417 9506 25469 9512
rect 25424 9466 25452 9506
rect 25240 9450 25452 9466
rect 25228 9444 25452 9450
rect 25280 9438 25452 9444
rect 25228 9386 25280 9392
rect 25136 8016 25188 8022
rect 25136 7958 25188 7964
rect 25148 7274 25176 7958
rect 25516 7324 25544 11047
rect 25700 9654 25728 12406
rect 25884 11830 25912 17478
rect 25976 15162 26004 21406
rect 26068 17610 26096 21626
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26056 17604 26108 17610
rect 26056 17546 26108 17552
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 25976 15065 26004 15098
rect 25962 15056 26018 15065
rect 25962 14991 26018 15000
rect 25964 14544 26016 14550
rect 25964 14486 26016 14492
rect 25976 12170 26004 14486
rect 26068 14006 26096 17274
rect 26160 15745 26188 21286
rect 26344 21128 26372 21830
rect 26528 21554 26556 21830
rect 26988 21690 27016 22102
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 26424 21140 26476 21146
rect 26344 21100 26424 21128
rect 26424 21082 26476 21088
rect 26988 21010 27016 21626
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26252 20602 26280 20810
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 20602 26464 20742
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26146 15736 26202 15745
rect 26146 15671 26202 15680
rect 26252 15620 26280 18906
rect 26422 18184 26478 18193
rect 26422 18119 26478 18128
rect 26160 15592 26280 15620
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 26160 13546 26188 15592
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26252 13734 26280 14554
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26160 13518 26280 13546
rect 26148 12640 26200 12646
rect 26148 12582 26200 12588
rect 26160 12238 26188 12582
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25872 11824 25924 11830
rect 25872 11766 25924 11772
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25792 10674 25820 11154
rect 25884 11150 25912 11290
rect 25976 11257 26004 11698
rect 26252 11286 26280 13518
rect 26344 11393 26372 14894
rect 26436 13530 26464 18119
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26424 13252 26476 13258
rect 26424 13194 26476 13200
rect 26436 12918 26464 13194
rect 26424 12912 26476 12918
rect 26424 12854 26476 12860
rect 26436 12238 26464 12854
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26330 11384 26386 11393
rect 26330 11319 26386 11328
rect 26240 11280 26292 11286
rect 25962 11248 26018 11257
rect 26240 11222 26292 11228
rect 26436 11218 26464 12174
rect 26528 11665 26556 19790
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26514 11656 26570 11665
rect 26514 11591 26570 11600
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 25962 11183 26018 11192
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 26436 11082 26464 11154
rect 26528 11150 26556 11494
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26332 11076 26384 11082
rect 26332 11018 26384 11024
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 26054 10976 26110 10985
rect 26054 10911 26110 10920
rect 26068 10826 26096 10911
rect 25976 10798 26096 10826
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25596 9648 25648 9654
rect 25688 9648 25740 9654
rect 25596 9590 25648 9596
rect 25686 9616 25688 9625
rect 25740 9616 25742 9625
rect 25608 9178 25636 9590
rect 25686 9551 25742 9560
rect 25700 9525 25728 9551
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25792 8548 25820 9386
rect 25872 8560 25924 8566
rect 25792 8520 25872 8548
rect 25872 8502 25924 8508
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25240 7296 25544 7324
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 24780 6582 24900 6610
rect 24780 6458 24808 6582
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24504 5494 24624 5522
rect 24504 4214 24532 5494
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 24688 4146 24716 4558
rect 24780 4146 24808 4966
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 24780 3058 24808 4082
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 24320 2378 24348 2790
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24136 870 24256 898
rect 24136 762 24164 870
rect 24228 800 24256 870
rect 24596 800 24624 2518
rect 24780 2514 24808 2994
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 24872 2446 24900 6394
rect 25148 6118 25176 7210
rect 25136 6112 25188 6118
rect 25134 6080 25136 6089
rect 25188 6080 25190 6089
rect 25134 6015 25190 6024
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24964 4554 24992 5170
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24964 800 24992 3878
rect 25240 3058 25268 7296
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 25332 5914 25360 6190
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25320 5296 25372 5302
rect 25320 5238 25372 5244
rect 25332 5098 25360 5238
rect 25320 5092 25372 5098
rect 25320 5034 25372 5040
rect 25332 4554 25360 5034
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4826 25452 4966
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25320 4548 25372 4554
rect 25320 4490 25372 4496
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25332 800 25360 2858
rect 25516 2446 25544 7142
rect 25608 6934 25636 7346
rect 25596 6928 25648 6934
rect 25596 6870 25648 6876
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25792 5817 25820 6054
rect 25778 5808 25834 5817
rect 25778 5743 25834 5752
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 25608 3194 25636 5170
rect 25700 4146 25728 5170
rect 25884 4146 25912 8502
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25686 3904 25742 3913
rect 25686 3839 25742 3848
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25700 800 25728 3839
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 25884 2990 25912 3538
rect 25976 3058 26004 10798
rect 26252 10266 26280 11018
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 26068 8566 26096 9386
rect 26252 8838 26280 9998
rect 26344 9654 26372 11018
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 26056 8560 26108 8566
rect 26056 8502 26108 8508
rect 26068 8294 26096 8502
rect 26252 8498 26280 8774
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26056 8288 26108 8294
rect 26056 8230 26108 8236
rect 26436 7818 26464 10202
rect 26620 9738 26648 18566
rect 26804 17746 26832 20878
rect 27172 18834 27200 22986
rect 27356 22778 27384 24704
rect 27896 24676 27948 24682
rect 27896 24618 27948 24624
rect 27712 24608 27764 24614
rect 27712 24550 27764 24556
rect 27724 24206 27752 24550
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27264 20534 27292 21082
rect 27448 20942 27476 24142
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27540 23050 27568 23190
rect 27528 23044 27580 23050
rect 27528 22986 27580 22992
rect 27540 22710 27568 22986
rect 27528 22704 27580 22710
rect 27724 22692 27752 24006
rect 27528 22646 27580 22652
rect 27632 22664 27752 22692
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27540 21729 27568 21830
rect 27526 21720 27582 21729
rect 27526 21655 27582 21664
rect 27540 21554 27568 21655
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27540 20942 27568 21490
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 27344 20324 27396 20330
rect 27344 20266 27396 20272
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27264 19514 27292 19722
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27172 18714 27200 18770
rect 27080 18686 27200 18714
rect 27080 18290 27108 18686
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 26792 17740 26844 17746
rect 26792 17682 26844 17688
rect 26804 16794 26832 17682
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26884 15632 26936 15638
rect 26884 15574 26936 15580
rect 26896 14550 26924 15574
rect 26988 15026 27016 16050
rect 27080 15706 27108 16934
rect 27068 15700 27120 15706
rect 27068 15642 27120 15648
rect 27066 15464 27122 15473
rect 27066 15399 27122 15408
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 26790 14376 26846 14385
rect 26790 14311 26846 14320
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26712 10985 26740 12038
rect 26698 10976 26754 10985
rect 26698 10911 26754 10920
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26528 9710 26648 9738
rect 26528 9489 26556 9710
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26514 9480 26570 9489
rect 26514 9415 26570 9424
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26424 7812 26476 7818
rect 26424 7754 26476 7760
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26068 5914 26096 6258
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 26068 4758 26096 4966
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 26056 4548 26108 4554
rect 26056 4490 26108 4496
rect 26068 3602 26096 4490
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 26160 3194 26188 7346
rect 26252 6866 26280 7754
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 26528 7410 26556 7686
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26252 3738 26280 6258
rect 26436 4146 26464 7346
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26528 4554 26556 6802
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26528 3670 26556 4014
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 26620 3534 26648 9590
rect 26712 6322 26740 9862
rect 26804 9586 26832 14311
rect 26884 14272 26936 14278
rect 26884 14214 26936 14220
rect 26896 13462 26924 14214
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26988 12850 27016 13670
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27080 12730 27108 15399
rect 26988 12702 27108 12730
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 26896 10849 26924 11154
rect 26882 10840 26938 10849
rect 26882 10775 26938 10784
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 26804 2774 26832 9318
rect 26896 8974 26924 9590
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 26896 7478 26924 8910
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 26896 6866 26924 7414
rect 26884 6860 26936 6866
rect 26884 6802 26936 6808
rect 26884 6724 26936 6730
rect 26884 6666 26936 6672
rect 26896 6458 26924 6666
rect 26988 6662 27016 12702
rect 27172 12374 27200 18566
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27264 12714 27292 13262
rect 27252 12708 27304 12714
rect 27252 12650 27304 12656
rect 27160 12368 27212 12374
rect 27160 12310 27212 12316
rect 27264 12238 27292 12650
rect 27356 12434 27384 20266
rect 27540 20058 27568 20878
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 27448 17066 27476 19450
rect 27632 19394 27660 22664
rect 27816 22642 27844 24346
rect 27908 24070 27936 24618
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 28000 23866 28028 24754
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 28184 23730 28212 25094
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 27804 22636 27856 22642
rect 27724 22596 27804 22624
rect 27724 22030 27752 22596
rect 27804 22578 27856 22584
rect 28080 22636 28132 22642
rect 28080 22578 28132 22584
rect 27804 22500 27856 22506
rect 27804 22442 27856 22448
rect 27896 22500 27948 22506
rect 27896 22442 27948 22448
rect 27816 22234 27844 22442
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27908 22030 27936 22442
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27896 22024 27948 22030
rect 27896 21966 27948 21972
rect 27988 21616 28040 21622
rect 28092 21604 28120 22578
rect 28184 22098 28212 23666
rect 28276 23526 28304 25842
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28368 23662 28396 24006
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 28040 21576 28120 21604
rect 27988 21558 28040 21564
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27724 21078 27752 21422
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27816 20992 27844 21286
rect 27896 21004 27948 21010
rect 27816 20964 27896 20992
rect 27816 20466 27844 20964
rect 27896 20946 27948 20952
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 28092 20330 28120 21576
rect 28080 20324 28132 20330
rect 28080 20266 28132 20272
rect 28184 20262 28212 22034
rect 28368 22030 28396 23598
rect 28460 22642 28488 24074
rect 28552 24070 28580 24754
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28644 23866 28672 25910
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 29368 25832 29420 25838
rect 29368 25774 29420 25780
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28632 23860 28684 23866
rect 28632 23802 28684 23808
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28262 21176 28318 21185
rect 28262 21111 28264 21120
rect 28316 21111 28318 21120
rect 28264 21082 28316 21088
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28080 19984 28132 19990
rect 28080 19926 28132 19932
rect 28092 19514 28120 19926
rect 28264 19780 28316 19786
rect 28264 19722 28316 19728
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27528 19372 27580 19378
rect 27632 19366 27936 19394
rect 27528 19314 27580 19320
rect 27540 18086 27568 19314
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27632 18970 27660 19246
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27712 18760 27764 18766
rect 27764 18720 27844 18748
rect 27712 18702 27764 18708
rect 27816 18290 27844 18720
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27620 18148 27672 18154
rect 27620 18090 27672 18096
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27436 17060 27488 17066
rect 27436 17002 27488 17008
rect 27448 16726 27476 17002
rect 27436 16720 27488 16726
rect 27436 16662 27488 16668
rect 27632 14414 27660 18090
rect 27816 17814 27844 18226
rect 27804 17808 27856 17814
rect 27804 17750 27856 17756
rect 27908 17218 27936 19366
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 28000 18290 28028 18770
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28092 18426 28120 18702
rect 28172 18692 28224 18698
rect 28172 18634 28224 18640
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28092 17882 28120 18362
rect 28184 18290 28212 18634
rect 28276 18358 28304 19722
rect 28368 18766 28396 21966
rect 28460 21554 28488 22170
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 19718 28488 20810
rect 28552 20602 28580 23598
rect 28644 23050 28672 23802
rect 29012 23798 29040 24550
rect 29000 23792 29052 23798
rect 29000 23734 29052 23740
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 28632 23044 28684 23050
rect 28684 23004 28764 23032
rect 28632 22986 28684 22992
rect 28736 21350 28764 23004
rect 28828 22778 28856 23530
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 29182 21584 29238 21593
rect 29182 21519 29184 21528
rect 29236 21519 29238 21528
rect 29184 21490 29236 21496
rect 28828 21457 29040 21468
rect 28814 21448 29054 21457
rect 28870 21440 28998 21448
rect 28814 21383 28870 21392
rect 28998 21383 29054 21392
rect 28724 21344 28776 21350
rect 29000 21344 29052 21350
rect 28776 21292 28948 21298
rect 28724 21286 28948 21292
rect 29000 21286 29052 21292
rect 28736 21270 28948 21286
rect 28814 21176 28870 21185
rect 28920 21146 28948 21270
rect 28814 21111 28870 21120
rect 28908 21140 28960 21146
rect 28828 21078 28856 21111
rect 28908 21082 28960 21088
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 29012 20942 29040 21286
rect 29288 21146 29316 23666
rect 29184 21140 29236 21146
rect 29184 21082 29236 21088
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29000 20936 29052 20942
rect 28632 20914 28684 20920
rect 29000 20878 29052 20884
rect 29104 20874 29132 20946
rect 29196 20874 29224 21082
rect 29380 21026 29408 25774
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 29840 24886 29868 25230
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 29828 24880 29880 24886
rect 29828 24822 29880 24828
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30288 24676 30340 24682
rect 30288 24618 30340 24624
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29840 24206 29868 24550
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29920 23792 29972 23798
rect 29920 23734 29972 23740
rect 29736 23180 29788 23186
rect 29736 23122 29788 23128
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 29656 22234 29684 22918
rect 29748 22778 29776 23122
rect 29736 22772 29788 22778
rect 29736 22714 29788 22720
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29644 22228 29696 22234
rect 29644 22170 29696 22176
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29564 21554 29592 22102
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 29656 21486 29684 21966
rect 29840 21962 29868 22714
rect 29932 22642 29960 23734
rect 30012 23112 30064 23118
rect 30010 23080 30012 23089
rect 30064 23080 30066 23089
rect 30010 23015 30066 23024
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22710 30144 22918
rect 30104 22704 30156 22710
rect 30024 22664 30104 22692
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 29920 22092 29972 22098
rect 29920 22034 29972 22040
rect 29932 22001 29960 22034
rect 29918 21992 29974 22001
rect 29828 21956 29880 21962
rect 29918 21927 29974 21936
rect 29828 21898 29880 21904
rect 30024 21554 30052 22664
rect 30300 22658 30328 24618
rect 30392 23254 30420 24754
rect 30484 23322 30512 25162
rect 30576 23798 30604 25842
rect 34796 25832 34848 25838
rect 34796 25774 34848 25780
rect 32864 25696 32916 25702
rect 32864 25638 32916 25644
rect 31668 25288 31720 25294
rect 31668 25230 31720 25236
rect 30748 25220 30800 25226
rect 30748 25162 30800 25168
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30576 23662 30604 23734
rect 30564 23656 30616 23662
rect 30564 23598 30616 23604
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30380 23248 30432 23254
rect 30380 23190 30432 23196
rect 30472 23112 30524 23118
rect 30472 23054 30524 23060
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30104 22646 30156 22652
rect 30208 22630 30328 22658
rect 30208 22522 30236 22630
rect 30116 22494 30236 22522
rect 30288 22568 30340 22574
rect 30288 22510 30340 22516
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 30116 21486 30144 22494
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 30208 21554 30236 22034
rect 30300 22030 30328 22510
rect 30392 22234 30420 22986
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30484 22094 30512 23054
rect 30564 23044 30616 23050
rect 30564 22986 30616 22992
rect 30576 22778 30604 22986
rect 30760 22778 30788 25162
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31220 24274 31248 25094
rect 31208 24268 31260 24274
rect 31208 24210 31260 24216
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 30852 22642 30880 24074
rect 30944 23118 30972 24142
rect 31312 24138 31340 25094
rect 31680 24206 31708 25230
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 31668 24200 31720 24206
rect 31668 24142 31720 24148
rect 31300 24132 31352 24138
rect 31300 24074 31352 24080
rect 32048 23798 32076 24686
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32036 23792 32088 23798
rect 32036 23734 32088 23740
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 31036 22642 31064 23122
rect 31404 23118 31432 23462
rect 31392 23112 31444 23118
rect 31206 23080 31262 23089
rect 31392 23054 31444 23060
rect 31206 23015 31208 23024
rect 31260 23015 31262 23024
rect 31208 22986 31260 22992
rect 31772 22642 31800 23666
rect 32048 22710 32076 23734
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32140 23526 32168 23666
rect 32128 23520 32180 23526
rect 32128 23462 32180 23468
rect 32324 23118 32352 24550
rect 32496 23792 32548 23798
rect 32692 23746 32720 24754
rect 32772 24404 32824 24410
rect 32772 24346 32824 24352
rect 32548 23740 32720 23746
rect 32496 23734 32720 23740
rect 32508 23718 32720 23734
rect 32784 23730 32812 24346
rect 32496 23180 32548 23186
rect 32496 23122 32548 23128
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32036 22704 32088 22710
rect 32036 22646 32088 22652
rect 30840 22636 30892 22642
rect 31021 22636 31073 22642
rect 30892 22596 30972 22624
rect 30840 22578 30892 22584
rect 30748 22568 30800 22574
rect 30748 22510 30800 22516
rect 30392 22066 30512 22094
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 29644 21480 29696 21486
rect 29644 21422 29696 21428
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 29920 21344 29972 21350
rect 29920 21286 29972 21292
rect 29932 21146 29960 21286
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 29288 20998 29408 21026
rect 28632 20856 28684 20862
rect 28724 20868 28776 20874
rect 28644 20602 28672 20856
rect 28724 20810 28776 20816
rect 29092 20868 29144 20874
rect 29092 20810 29144 20816
rect 29184 20868 29236 20874
rect 29184 20810 29236 20816
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 28736 20398 28764 20810
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28448 19712 28500 19718
rect 28448 19654 28500 19660
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28184 17338 28212 18226
rect 28264 18216 28316 18222
rect 28368 18204 28396 18702
rect 28316 18176 28396 18204
rect 28264 18158 28316 18164
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 27908 17190 28304 17218
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27724 16114 27752 17002
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27724 15162 27752 16050
rect 27816 15609 27844 16526
rect 27908 16046 27936 17070
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28184 16114 28212 16390
rect 27988 16108 28040 16114
rect 28172 16108 28224 16114
rect 28040 16068 28120 16096
rect 27988 16050 28040 16056
rect 27896 16040 27948 16046
rect 27896 15982 27948 15988
rect 27802 15600 27858 15609
rect 27802 15535 27858 15544
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27724 14346 27752 15098
rect 27816 14482 27844 15535
rect 27908 15434 27936 15982
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27908 15094 27936 15370
rect 27896 15088 27948 15094
rect 27896 15030 27948 15036
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 13938 27476 14214
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27712 13252 27764 13258
rect 27712 13194 27764 13200
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27356 12406 27476 12434
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 27068 10464 27120 10470
rect 27068 10406 27120 10412
rect 27080 9654 27108 10406
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27066 8936 27122 8945
rect 27066 8871 27068 8880
rect 27120 8871 27122 8880
rect 27068 8842 27120 8848
rect 27172 8498 27200 11222
rect 27264 10130 27292 12174
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27356 10198 27384 11222
rect 27448 10962 27476 12406
rect 27540 11762 27568 13126
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27632 12306 27660 12786
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27540 11121 27568 11698
rect 27526 11112 27582 11121
rect 27526 11047 27582 11056
rect 27448 10934 27568 10962
rect 27540 10538 27568 10934
rect 27632 10674 27660 12242
rect 27724 11830 27752 13194
rect 27908 12646 27936 13194
rect 27896 12640 27948 12646
rect 27896 12582 27948 12588
rect 28000 12434 28028 14962
rect 27908 12406 28028 12434
rect 27712 11824 27764 11830
rect 27712 11766 27764 11772
rect 27724 11150 27752 11766
rect 27712 11144 27764 11150
rect 27712 11086 27764 11092
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27344 10192 27396 10198
rect 27344 10134 27396 10140
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 27264 9568 27292 10066
rect 27344 9580 27396 9586
rect 27264 9540 27344 9568
rect 27264 8974 27292 9540
rect 27344 9522 27396 9528
rect 27540 9081 27568 10474
rect 27632 9518 27660 10610
rect 27724 10062 27752 11086
rect 27816 10985 27844 11086
rect 27802 10976 27858 10985
rect 27802 10911 27858 10920
rect 27908 10146 27936 12406
rect 27986 12336 28042 12345
rect 27986 12271 28042 12280
rect 27816 10118 27936 10146
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27710 9480 27766 9489
rect 27710 9415 27766 9424
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27632 9217 27660 9318
rect 27618 9208 27674 9217
rect 27618 9143 27674 9152
rect 27526 9072 27582 9081
rect 27436 9036 27488 9042
rect 27526 9007 27582 9016
rect 27436 8978 27488 8984
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27344 8832 27396 8838
rect 27344 8774 27396 8780
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27080 7818 27108 8366
rect 27068 7812 27120 7818
rect 27068 7754 27120 7760
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26882 5672 26938 5681
rect 26882 5607 26884 5616
rect 26936 5607 26938 5616
rect 26976 5636 27028 5642
rect 26884 5578 26936 5584
rect 26976 5578 27028 5584
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 26896 4622 26924 4966
rect 26884 4616 26936 4622
rect 26884 4558 26936 4564
rect 26896 4146 26924 4558
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26896 3534 26924 3878
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 26988 3058 27016 5578
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 27080 4826 27108 4966
rect 27068 4820 27120 4826
rect 27068 4762 27120 4768
rect 27172 4622 27200 8434
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26252 2746 26832 2774
rect 26252 2378 26280 2746
rect 27080 2514 27108 4490
rect 27264 3602 27292 8026
rect 27356 4146 27384 8774
rect 27448 7886 27476 8978
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27540 8430 27568 8910
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27540 7834 27568 8026
rect 27540 7806 27660 7834
rect 27528 7744 27580 7750
rect 27434 7712 27490 7721
rect 27528 7686 27580 7692
rect 27434 7647 27490 7656
rect 27448 6798 27476 7647
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27434 5808 27490 5817
rect 27434 5743 27436 5752
rect 27488 5743 27490 5752
rect 27436 5714 27488 5720
rect 27540 5710 27568 7686
rect 27632 7478 27660 7806
rect 27620 7472 27672 7478
rect 27620 7414 27672 7420
rect 27724 6882 27752 9415
rect 27816 7154 27844 10118
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27908 9722 27936 9930
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27894 9344 27950 9353
rect 27894 9279 27950 9288
rect 27908 8566 27936 9279
rect 27896 8560 27948 8566
rect 27896 8502 27948 8508
rect 28000 7313 28028 12271
rect 28092 11540 28120 16068
rect 28172 16050 28224 16056
rect 28276 15994 28304 17190
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28368 16114 28396 16458
rect 28460 16114 28488 16934
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28184 15966 28304 15994
rect 28184 12345 28212 15966
rect 28368 15570 28396 16050
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28276 14618 28304 15438
rect 28368 15026 28396 15506
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28460 14498 28488 16050
rect 28552 15978 28580 20334
rect 28724 20256 28776 20262
rect 28724 20198 28776 20204
rect 28630 19272 28686 19281
rect 28630 19207 28632 19216
rect 28684 19207 28686 19216
rect 28632 19178 28684 19184
rect 28736 18766 28764 20198
rect 28816 19780 28868 19786
rect 28816 19722 28868 19728
rect 28828 19446 28856 19722
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28736 18290 28764 18702
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28736 17134 28764 18226
rect 28920 18154 28948 20538
rect 29288 19334 29316 20998
rect 29552 20800 29604 20806
rect 29552 20742 29604 20748
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29564 19854 29592 20742
rect 29840 20602 29868 20742
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29104 19306 29316 19334
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29104 18834 29132 19306
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28724 15972 28776 15978
rect 28724 15914 28776 15920
rect 28276 14470 28488 14498
rect 28540 14476 28592 14482
rect 28170 12336 28226 12345
rect 28170 12271 28226 12280
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28184 11898 28212 12174
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28276 11694 28304 14470
rect 28540 14418 28592 14424
rect 28356 14272 28408 14278
rect 28356 14214 28408 14220
rect 28264 11688 28316 11694
rect 28264 11630 28316 11636
rect 28092 11512 28304 11540
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 28092 8362 28120 11018
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28184 9450 28212 9930
rect 28172 9444 28224 9450
rect 28172 9386 28224 9392
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 28184 8673 28212 8774
rect 28170 8664 28226 8673
rect 28170 8599 28226 8608
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 28184 7818 28212 8230
rect 28172 7812 28224 7818
rect 28172 7754 28224 7760
rect 28184 7410 28212 7754
rect 28276 7449 28304 11512
rect 28368 8974 28396 14214
rect 28552 13870 28580 14418
rect 28736 14006 28764 15914
rect 28920 15910 28948 18090
rect 29012 17592 29040 18566
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29104 17762 29132 18226
rect 29196 17882 29224 19110
rect 29276 18760 29328 18766
rect 29276 18702 29328 18708
rect 29288 18222 29316 18702
rect 29380 18426 29408 19314
rect 29460 18896 29512 18902
rect 29460 18838 29512 18844
rect 29368 18420 29420 18426
rect 29368 18362 29420 18368
rect 29276 18216 29328 18222
rect 29276 18158 29328 18164
rect 29184 17876 29236 17882
rect 29184 17818 29236 17824
rect 29104 17734 29224 17762
rect 29092 17604 29144 17610
rect 29012 17564 29092 17592
rect 29012 17202 29040 17564
rect 29092 17546 29144 17552
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29196 17066 29224 17734
rect 29288 17066 29316 18158
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29380 17678 29408 18022
rect 29368 17672 29420 17678
rect 29368 17614 29420 17620
rect 29472 17542 29500 18838
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 29564 17338 29592 19314
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29656 18970 29684 19246
rect 29748 19174 29776 20402
rect 29932 20330 29960 21082
rect 29920 20324 29972 20330
rect 29920 20266 29972 20272
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29644 18964 29696 18970
rect 29644 18906 29696 18912
rect 29656 17882 29684 18906
rect 29748 18290 29776 19110
rect 30116 18698 30144 21422
rect 30208 21078 30236 21490
rect 30300 21350 30328 21966
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 30196 21072 30248 21078
rect 30196 21014 30248 21020
rect 30288 20460 30340 20466
rect 30392 20448 30420 22066
rect 30564 21480 30616 21486
rect 30760 21457 30788 22510
rect 30564 21422 30616 21428
rect 30746 21448 30802 21457
rect 30576 20942 30604 21422
rect 30746 21383 30802 21392
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30340 20420 30420 20448
rect 30288 20402 30340 20408
rect 30288 20324 30340 20330
rect 30288 20266 30340 20272
rect 30300 18970 30328 20266
rect 30392 19446 30420 20420
rect 30472 20392 30524 20398
rect 30472 20334 30524 20340
rect 30484 19854 30512 20334
rect 30576 20058 30604 20878
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 30380 19236 30432 19242
rect 30380 19178 30432 19184
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30196 18760 30248 18766
rect 30248 18720 30328 18748
rect 30196 18702 30248 18708
rect 30104 18692 30156 18698
rect 30104 18634 30156 18640
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29644 17876 29696 17882
rect 29644 17818 29696 17824
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29184 17060 29236 17066
rect 29184 17002 29236 17008
rect 29276 17060 29328 17066
rect 29276 17002 29328 17008
rect 29196 16726 29224 17002
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29184 16720 29236 16726
rect 29184 16662 29236 16668
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28828 15502 28856 15846
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28816 14884 28868 14890
rect 28816 14826 28868 14832
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 28644 12850 28672 13942
rect 28828 13326 28856 14826
rect 28920 14414 28948 15846
rect 29564 15570 29592 16730
rect 29748 16658 29776 18226
rect 30116 18222 30144 18634
rect 30300 18290 30328 18720
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 30300 16250 30328 18226
rect 30392 16590 30420 19178
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30484 17814 30512 18702
rect 30576 18426 30604 18702
rect 30668 18426 30696 19790
rect 30852 19378 30880 20742
rect 30944 19854 30972 22596
rect 31021 22578 31073 22584
rect 31116 22636 31168 22642
rect 31760 22636 31812 22642
rect 31168 22596 31248 22624
rect 31116 22578 31168 22584
rect 31220 21690 31248 22596
rect 31760 22578 31812 22584
rect 32140 22030 32168 23054
rect 32416 22778 32444 23054
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 31312 21554 31340 21966
rect 32324 21554 32352 22578
rect 32508 22166 32536 23122
rect 32692 22642 32720 23718
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 32876 23594 32904 25638
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 32956 24132 33008 24138
rect 32956 24074 33008 24080
rect 33048 24132 33100 24138
rect 33100 24092 33180 24120
rect 33048 24074 33100 24080
rect 32968 23866 32996 24074
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 32956 23724 33008 23730
rect 32956 23666 33008 23672
rect 32772 23588 32824 23594
rect 32772 23530 32824 23536
rect 32864 23588 32916 23594
rect 32864 23530 32916 23536
rect 32784 23474 32812 23530
rect 32968 23474 32996 23666
rect 32784 23446 32996 23474
rect 32956 23180 33008 23186
rect 32956 23122 33008 23128
rect 32864 22976 32916 22982
rect 32864 22918 32916 22924
rect 32876 22710 32904 22918
rect 32772 22704 32824 22710
rect 32772 22646 32824 22652
rect 32864 22704 32916 22710
rect 32864 22646 32916 22652
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32692 22250 32720 22578
rect 32600 22222 32720 22250
rect 32496 22160 32548 22166
rect 32496 22102 32548 22108
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 31300 21548 31352 21554
rect 31300 21490 31352 21496
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32312 21412 32364 21418
rect 32312 21354 32364 21360
rect 32324 21146 32352 21354
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32416 21010 32444 21490
rect 32508 21146 32536 21966
rect 32496 21140 32548 21146
rect 32496 21082 32548 21088
rect 32404 21004 32456 21010
rect 32404 20946 32456 20952
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 31404 19922 31432 20402
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 30932 19440 30984 19446
rect 30932 19382 30984 19388
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30564 18420 30616 18426
rect 30564 18362 30616 18368
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30472 17808 30524 17814
rect 30472 17750 30524 17756
rect 30852 17338 30880 19314
rect 30944 18290 30972 19382
rect 31036 18358 31064 19790
rect 32324 19514 32352 20878
rect 32600 20602 32628 22222
rect 32680 22092 32732 22098
rect 32680 22034 32732 22040
rect 32692 21690 32720 22034
rect 32680 21684 32732 21690
rect 32680 21626 32732 21632
rect 32784 21078 32812 22646
rect 32864 21548 32916 21554
rect 32864 21490 32916 21496
rect 32876 21078 32904 21490
rect 32772 21072 32824 21078
rect 32772 21014 32824 21020
rect 32864 21072 32916 21078
rect 32864 21014 32916 21020
rect 32784 20806 32812 21014
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32772 20596 32824 20602
rect 32772 20538 32824 20544
rect 32588 19848 32640 19854
rect 32588 19790 32640 19796
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32220 18964 32272 18970
rect 32220 18906 32272 18912
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 31024 18352 31076 18358
rect 31024 18294 31076 18300
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30944 18154 30972 18226
rect 30932 18148 30984 18154
rect 30932 18090 30984 18096
rect 30944 17678 30972 18090
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 31036 17610 31064 18294
rect 31392 18148 31444 18154
rect 31392 18090 31444 18096
rect 31404 17678 31432 18090
rect 31760 18080 31812 18086
rect 31760 18022 31812 18028
rect 31772 17746 31800 18022
rect 32048 17814 32076 18702
rect 32036 17808 32088 17814
rect 32036 17750 32088 17756
rect 32232 17746 32260 18906
rect 32416 18358 32444 19314
rect 32600 19122 32628 19790
rect 32600 19094 32720 19122
rect 32692 18714 32720 19094
rect 32784 18902 32812 20538
rect 32876 20058 32904 21014
rect 32968 20602 32996 23122
rect 33152 22642 33180 24092
rect 33416 23860 33468 23866
rect 33244 23820 33416 23848
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33244 22574 33272 23820
rect 33416 23802 33468 23808
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 33796 23594 33824 23666
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 33784 23588 33836 23594
rect 33784 23530 33836 23536
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33232 22568 33284 22574
rect 33232 22510 33284 22516
rect 33336 22438 33364 23054
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 22522 33456 22578
rect 33428 22494 33548 22522
rect 33324 22432 33376 22438
rect 33324 22374 33376 22380
rect 33336 22234 33364 22374
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 32956 20596 33008 20602
rect 32956 20538 33008 20544
rect 32864 20052 32916 20058
rect 32864 19994 32916 20000
rect 33060 19854 33088 21966
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 33152 21622 33180 21830
rect 33140 21616 33192 21622
rect 33140 21558 33192 21564
rect 33336 21010 33364 22034
rect 33520 21486 33548 22494
rect 33600 21956 33652 21962
rect 33600 21898 33652 21904
rect 33612 21690 33640 21898
rect 33600 21684 33652 21690
rect 33600 21626 33652 21632
rect 33876 21616 33928 21622
rect 33876 21558 33928 21564
rect 33508 21480 33560 21486
rect 33508 21422 33560 21428
rect 33324 21004 33376 21010
rect 33324 20946 33376 20952
rect 33416 20800 33468 20806
rect 33416 20742 33468 20748
rect 33428 20534 33456 20742
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33520 20466 33548 21422
rect 33888 20942 33916 21558
rect 33876 20936 33928 20942
rect 33876 20878 33928 20884
rect 33324 20460 33376 20466
rect 33324 20402 33376 20408
rect 33508 20460 33560 20466
rect 33508 20402 33560 20408
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 32956 19712 33008 19718
rect 32956 19654 33008 19660
rect 32968 19514 32996 19654
rect 32956 19508 33008 19514
rect 32956 19450 33008 19456
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 32772 18896 32824 18902
rect 32772 18838 32824 18844
rect 32692 18686 32812 18714
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32496 18420 32548 18426
rect 32496 18362 32548 18368
rect 32404 18352 32456 18358
rect 32404 18294 32456 18300
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31036 17338 31064 17546
rect 32232 17542 32260 17682
rect 32416 17678 32444 18294
rect 32508 17678 32536 18362
rect 32600 18290 32628 18566
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 32220 17536 32272 17542
rect 32220 17478 32272 17484
rect 30472 17332 30524 17338
rect 30472 17274 30524 17280
rect 30840 17332 30892 17338
rect 30840 17274 30892 17280
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 30484 16794 30512 17274
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31668 17196 31720 17202
rect 31668 17138 31720 17144
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 30840 17060 30892 17066
rect 30840 17002 30892 17008
rect 30472 16788 30524 16794
rect 30472 16730 30524 16736
rect 30852 16726 30880 17002
rect 30840 16720 30892 16726
rect 30840 16662 30892 16668
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30472 16516 30524 16522
rect 30472 16458 30524 16464
rect 30288 16244 30340 16250
rect 30288 16186 30340 16192
rect 30484 15978 30512 16458
rect 31036 16046 31064 17138
rect 31680 16590 31708 17138
rect 32232 16998 32260 17138
rect 32220 16992 32272 16998
rect 32220 16934 32272 16940
rect 32232 16658 32260 16934
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 31668 16584 31720 16590
rect 31668 16526 31720 16532
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 30656 16040 30708 16046
rect 30656 15982 30708 15988
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 30472 15972 30524 15978
rect 30472 15914 30524 15920
rect 30484 15706 30512 15914
rect 30472 15700 30524 15706
rect 30472 15642 30524 15648
rect 29276 15564 29328 15570
rect 29276 15506 29328 15512
rect 29552 15564 29604 15570
rect 29552 15506 29604 15512
rect 29288 15026 29316 15506
rect 30668 15502 30696 15982
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 29368 15360 29420 15366
rect 29368 15302 29420 15308
rect 29380 15026 29408 15302
rect 30668 15162 30696 15438
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 31220 15094 31248 16050
rect 31680 16046 31708 16526
rect 32128 16448 32180 16454
rect 32128 16390 32180 16396
rect 32140 16114 32168 16390
rect 32416 16250 32444 17614
rect 32600 17338 32628 18226
rect 32784 17678 32812 18686
rect 32876 18222 32904 19382
rect 33152 19310 33180 19858
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33336 18970 33364 20402
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33232 18828 33284 18834
rect 33232 18770 33284 18776
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 32956 18692 33008 18698
rect 32956 18634 33008 18640
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32772 17672 32824 17678
rect 32772 17614 32824 17620
rect 32876 17542 32904 18158
rect 32968 18086 32996 18634
rect 33152 18086 33180 18702
rect 33244 18290 33272 18770
rect 33324 18624 33376 18630
rect 33324 18566 33376 18572
rect 33232 18284 33284 18290
rect 33232 18226 33284 18232
rect 32956 18080 33008 18086
rect 32956 18022 33008 18028
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 32864 17536 32916 17542
rect 32864 17478 32916 17484
rect 32588 17332 32640 17338
rect 32588 17274 32640 17280
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 32956 16584 33008 16590
rect 33060 16574 33088 16934
rect 33152 16658 33180 18022
rect 33336 17882 33364 18566
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 33428 17746 33456 19790
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33796 19514 33824 19722
rect 33784 19508 33836 19514
rect 33784 19450 33836 19456
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33612 18290 33640 18362
rect 33692 18352 33744 18358
rect 33876 18352 33928 18358
rect 33744 18312 33876 18340
rect 33692 18294 33744 18300
rect 33876 18294 33928 18300
rect 34164 18290 34192 23598
rect 34440 23594 34468 23666
rect 34428 23588 34480 23594
rect 34428 23530 34480 23536
rect 34716 23118 34744 24346
rect 34808 23322 34836 25774
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 34704 23112 34756 23118
rect 34704 23054 34756 23060
rect 34716 22030 34744 23054
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34808 21554 34836 22034
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 20602 34836 21490
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34796 20596 34848 20602
rect 34796 20538 34848 20544
rect 34808 19446 34836 20538
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35360 19990 35388 46990
rect 35622 21992 35678 22001
rect 35622 21927 35678 21936
rect 35636 21486 35664 21927
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35348 19984 35400 19990
rect 35348 19926 35400 19932
rect 34796 19440 34848 19446
rect 34796 19382 34848 19388
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34164 18086 34192 18226
rect 34152 18080 34204 18086
rect 34152 18022 34204 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 33416 17740 33468 17746
rect 33416 17682 33468 17688
rect 33428 17610 33456 17682
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33416 17604 33468 17610
rect 33416 17546 33468 17552
rect 33324 17196 33376 17202
rect 33324 17138 33376 17144
rect 33140 16652 33192 16658
rect 33140 16594 33192 16600
rect 33008 16546 33088 16574
rect 32956 16526 33008 16532
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32128 16108 32180 16114
rect 32128 16050 32180 16056
rect 31668 16040 31720 16046
rect 31668 15982 31720 15988
rect 31680 15570 31708 15982
rect 32968 15910 32996 16526
rect 33336 16250 33364 17138
rect 33428 16794 33456 17546
rect 33612 17338 33640 17614
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33324 16244 33376 16250
rect 33324 16186 33376 16192
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 31668 15564 31720 15570
rect 31668 15506 31720 15512
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 29276 15020 29328 15026
rect 29276 14962 29328 14968
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 28908 14408 28960 14414
rect 28908 14350 28960 14356
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 28816 13320 28868 13326
rect 28816 13262 28868 13268
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28460 11354 28488 12106
rect 28644 11762 28672 12786
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28736 10713 28764 11086
rect 28722 10704 28778 10713
rect 28722 10639 28778 10648
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10130 28764 10542
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28460 8498 28488 9454
rect 28538 8936 28594 8945
rect 28538 8871 28594 8880
rect 28552 8634 28580 8871
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28460 7936 28488 8434
rect 28828 8378 28856 12582
rect 28920 11898 28948 13126
rect 29012 12918 29040 13670
rect 29104 13462 29132 14282
rect 29196 14074 29224 14894
rect 29288 14482 29316 14962
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29656 14414 29684 14758
rect 31220 14618 31248 15030
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 31208 14612 31260 14618
rect 31208 14554 31260 14560
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29196 13530 29224 13874
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29092 13456 29144 13462
rect 29092 13398 29144 13404
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 29552 12096 29604 12102
rect 29552 12038 29604 12044
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 29564 11830 29592 12038
rect 29552 11824 29604 11830
rect 29552 11766 29604 11772
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 29092 11348 29144 11354
rect 29092 11290 29144 11296
rect 31484 11348 31536 11354
rect 31484 11290 31536 11296
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28920 10810 28948 10950
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9042 29040 9998
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 28920 8566 28948 8978
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 28736 8350 28856 8378
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28540 7948 28592 7954
rect 28460 7908 28540 7936
rect 28540 7890 28592 7896
rect 28540 7744 28592 7750
rect 28644 7732 28672 7958
rect 28592 7704 28672 7732
rect 28540 7686 28592 7692
rect 28262 7440 28318 7449
rect 28172 7404 28224 7410
rect 28262 7375 28318 7384
rect 28172 7346 28224 7352
rect 27986 7304 28042 7313
rect 27986 7239 28042 7248
rect 27816 7126 28028 7154
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27632 6866 27844 6882
rect 27632 6860 27856 6866
rect 27632 6854 27804 6860
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27448 4282 27476 5102
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27632 3466 27660 6854
rect 27804 6802 27856 6808
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 5914 27844 6666
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27724 5302 27752 5646
rect 27712 5296 27764 5302
rect 27712 5238 27764 5244
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27252 3392 27304 3398
rect 27252 3334 27304 3340
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 26068 800 26096 2246
rect 26436 800 26464 2382
rect 26884 2372 26936 2378
rect 26884 2314 26936 2320
rect 26896 800 26924 2314
rect 27264 800 27292 3334
rect 27724 2922 27752 3538
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27816 3058 27844 3470
rect 27908 3398 27936 6938
rect 28000 5953 28028 7126
rect 28184 6798 28212 7346
rect 28356 7268 28408 7274
rect 28356 7210 28408 7216
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 27986 5944 28042 5953
rect 27986 5879 28042 5888
rect 28092 5681 28120 6190
rect 28172 6112 28224 6118
rect 28172 6054 28224 6060
rect 28264 6112 28316 6118
rect 28264 6054 28316 6060
rect 28078 5672 28134 5681
rect 28078 5607 28134 5616
rect 28184 4185 28212 6054
rect 28170 4176 28226 4185
rect 28170 4111 28172 4120
rect 28224 4111 28226 4120
rect 28172 4082 28224 4088
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28184 3126 28212 4082
rect 28276 3534 28304 6054
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 28172 3120 28224 3126
rect 28172 3062 28224 3068
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 27632 800 27660 2790
rect 28368 2446 28396 7210
rect 28552 6798 28580 7686
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28540 6792 28592 6798
rect 28540 6734 28592 6740
rect 28552 5302 28580 6734
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 28644 5216 28672 7482
rect 28736 6118 28764 8350
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28828 6866 28856 8230
rect 29012 7886 29040 8842
rect 29104 8809 29132 11290
rect 31496 11257 31524 11290
rect 31482 11248 31538 11257
rect 31482 11183 31538 11192
rect 29552 11144 29604 11150
rect 29828 11144 29880 11150
rect 29604 11104 29828 11132
rect 29552 11086 29604 11092
rect 29828 11086 29880 11092
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 29564 10674 29592 10950
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 30472 10668 30524 10674
rect 30472 10610 30524 10616
rect 30012 10124 30064 10130
rect 30012 10066 30064 10072
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29564 9897 29592 9998
rect 29550 9888 29606 9897
rect 29550 9823 29606 9832
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29090 8800 29146 8809
rect 29090 8735 29146 8744
rect 29196 8090 29224 8978
rect 29368 8968 29420 8974
rect 29656 8922 29684 9454
rect 29840 9178 29868 9998
rect 29828 9172 29880 9178
rect 29828 9114 29880 9120
rect 29368 8910 29420 8916
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29000 7880 29052 7886
rect 29000 7822 29052 7828
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28920 7478 28948 7686
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 29196 7410 29224 7890
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29196 6866 29224 7346
rect 28816 6860 28868 6866
rect 28816 6802 28868 6808
rect 29184 6860 29236 6866
rect 29184 6802 29236 6808
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 29288 6390 29316 6598
rect 29380 6474 29408 8910
rect 29472 8894 29684 8922
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29472 8838 29500 8894
rect 29460 8832 29512 8838
rect 29460 8774 29512 8780
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29564 7206 29592 7686
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29380 6446 29592 6474
rect 29276 6384 29328 6390
rect 29276 6326 29328 6332
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28816 5704 28868 5710
rect 29000 5704 29052 5710
rect 28868 5664 28948 5692
rect 28816 5646 28868 5652
rect 28920 5574 28948 5664
rect 29000 5646 29052 5652
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 28736 5352 28764 5510
rect 28908 5364 28960 5370
rect 28736 5324 28908 5352
rect 28908 5306 28960 5312
rect 28644 5188 28764 5216
rect 28632 5092 28684 5098
rect 28632 5034 28684 5040
rect 28540 4480 28592 4486
rect 28644 4468 28672 5034
rect 28592 4440 28672 4468
rect 28540 4422 28592 4428
rect 28644 3534 28672 4440
rect 28736 3602 28764 5188
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28828 4826 28856 4966
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28920 4554 28948 5306
rect 28908 4548 28960 4554
rect 28908 4490 28960 4496
rect 28814 4176 28870 4185
rect 28814 4111 28816 4120
rect 28868 4111 28870 4120
rect 28816 4082 28868 4088
rect 28920 3670 28948 4490
rect 29012 3738 29040 5646
rect 29288 5302 29316 6326
rect 29380 5846 29408 6326
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29472 5914 29500 6054
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29368 5840 29420 5846
rect 29368 5782 29420 5788
rect 29380 5710 29408 5782
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29276 5296 29328 5302
rect 29276 5238 29328 5244
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 29104 4214 29132 4558
rect 29564 4298 29592 6446
rect 29656 6322 29684 8774
rect 29840 8430 29868 8774
rect 29828 8424 29880 8430
rect 29828 8366 29880 8372
rect 29736 8356 29788 8362
rect 29736 8298 29788 8304
rect 29748 6458 29776 8298
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29748 5234 29776 6054
rect 29840 5642 29868 7142
rect 29932 6769 29960 8910
rect 29918 6760 29974 6769
rect 29918 6695 29974 6704
rect 30024 5846 30052 10066
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30116 6118 30144 9590
rect 30208 8498 30236 9862
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30208 6798 30236 8230
rect 30300 7478 30328 9862
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30392 9178 30420 9522
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30288 7472 30340 7478
rect 30288 7414 30340 7420
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30012 5840 30064 5846
rect 30012 5782 30064 5788
rect 30300 5778 30328 6258
rect 30392 5846 30420 8910
rect 30484 8634 30512 10610
rect 30852 10470 30880 10950
rect 31576 10668 31628 10674
rect 31576 10610 31628 10616
rect 31300 10532 31352 10538
rect 31300 10474 31352 10480
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 30932 9988 30984 9994
rect 30932 9930 30984 9936
rect 30746 9888 30802 9897
rect 30746 9823 30802 9832
rect 30760 9654 30788 9823
rect 30748 9648 30800 9654
rect 30748 9590 30800 9596
rect 30564 9580 30616 9586
rect 30564 9522 30616 9528
rect 30576 9489 30604 9522
rect 30562 9480 30618 9489
rect 30562 9415 30618 9424
rect 30654 9072 30710 9081
rect 30654 9007 30710 9016
rect 30668 8634 30696 9007
rect 30472 8628 30524 8634
rect 30656 8628 30708 8634
rect 30524 8588 30604 8616
rect 30472 8570 30524 8576
rect 30576 6866 30604 8588
rect 30656 8570 30708 8576
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30668 7818 30696 8434
rect 30656 7812 30708 7818
rect 30656 7754 30708 7760
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30760 6730 30788 9590
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30748 6724 30800 6730
rect 30748 6666 30800 6672
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29736 5228 29788 5234
rect 29736 5170 29788 5176
rect 29840 4690 29868 5578
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 29920 5296 29972 5302
rect 29920 5238 29972 5244
rect 29828 4684 29880 4690
rect 29828 4626 29880 4632
rect 29828 4548 29880 4554
rect 29828 4490 29880 4496
rect 29472 4282 29592 4298
rect 29460 4276 29592 4282
rect 29512 4270 29592 4276
rect 29460 4218 29512 4224
rect 29840 4214 29868 4490
rect 29932 4486 29960 5238
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 29920 4480 29972 4486
rect 29920 4422 29972 4428
rect 29932 4282 29960 4422
rect 30208 4282 30236 4966
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 29920 4276 29972 4282
rect 29920 4218 29972 4224
rect 30196 4276 30248 4282
rect 30196 4218 30248 4224
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29828 4208 29880 4214
rect 29828 4150 29880 4156
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28724 3596 28776 3602
rect 28724 3538 28776 3544
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28460 3058 28488 3334
rect 28920 3058 28948 3606
rect 29840 3602 29868 4150
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 30024 3602 30052 4082
rect 29828 3596 29880 3602
rect 29828 3538 29880 3544
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 30208 3534 30236 4218
rect 30300 4146 30328 4422
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 3194 29132 3334
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28736 2825 28764 2926
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 29000 2848 29052 2854
rect 28722 2816 28778 2825
rect 29000 2790 29052 2796
rect 28722 2751 28778 2760
rect 29012 2650 29040 2790
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28356 1420 28408 1426
rect 28356 1362 28408 1368
rect 28368 800 28396 1362
rect 29104 800 29132 2858
rect 29748 2854 29776 3470
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 29828 2304 29880 2310
rect 29828 2246 29880 2252
rect 29840 1426 29868 2246
rect 29828 1420 29880 1426
rect 29828 1362 29880 1368
rect 30024 1306 30052 3130
rect 30392 2446 30420 5510
rect 30484 5370 30512 6258
rect 30852 6254 30880 9318
rect 30944 8974 30972 9930
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 31036 6610 31064 10406
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31128 9110 31156 9318
rect 31116 9104 31168 9110
rect 31116 9046 31168 9052
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31128 8090 31156 8910
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31116 7472 31168 7478
rect 31116 7414 31168 7420
rect 30944 6582 31064 6610
rect 30840 6248 30892 6254
rect 30840 6190 30892 6196
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30760 4826 30788 5646
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 30564 2576 30616 2582
rect 30564 2518 30616 2524
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 29840 1278 30052 1306
rect 29840 800 29868 1278
rect 30576 800 30604 2518
rect 30852 2514 30880 5170
rect 30840 2508 30892 2514
rect 30840 2450 30892 2456
rect 30944 2106 30972 6582
rect 31128 6390 31156 7414
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31116 6384 31168 6390
rect 31116 6326 31168 6332
rect 31220 6254 31248 7142
rect 31312 6905 31340 10474
rect 31392 10056 31444 10062
rect 31392 9998 31444 10004
rect 31298 6896 31354 6905
rect 31298 6831 31354 6840
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 31208 6248 31260 6254
rect 31208 6190 31260 6196
rect 31024 6112 31076 6118
rect 31024 6054 31076 6060
rect 31036 2446 31064 6054
rect 31220 5914 31248 6190
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31312 5642 31340 6598
rect 31300 5636 31352 5642
rect 31300 5578 31352 5584
rect 31404 4706 31432 9998
rect 31484 9920 31536 9926
rect 31484 9862 31536 9868
rect 31496 9450 31524 9862
rect 31484 9444 31536 9450
rect 31484 9386 31536 9392
rect 31588 7002 31616 10610
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 31944 9580 31996 9586
rect 31944 9522 31996 9528
rect 33600 9580 33652 9586
rect 33600 9522 33652 9528
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31576 6996 31628 7002
rect 31576 6938 31628 6944
rect 31772 6905 31800 9318
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31482 6896 31538 6905
rect 31482 6831 31538 6840
rect 31758 6896 31814 6905
rect 31758 6831 31814 6840
rect 31128 4678 31432 4706
rect 31128 3466 31156 4678
rect 31300 4548 31352 4554
rect 31300 4490 31352 4496
rect 31312 3942 31340 4490
rect 31496 4026 31524 6831
rect 31864 6746 31892 8298
rect 31956 7585 31984 9522
rect 32496 9376 32548 9382
rect 32496 9318 32548 9324
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 32220 9104 32272 9110
rect 32220 9046 32272 9052
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 32140 8022 32168 8774
rect 32128 8016 32180 8022
rect 32128 7958 32180 7964
rect 32036 7812 32088 7818
rect 32036 7754 32088 7760
rect 31942 7576 31998 7585
rect 31942 7511 31998 7520
rect 31944 7336 31996 7342
rect 31944 7278 31996 7284
rect 31956 6798 31984 7278
rect 31668 6724 31720 6730
rect 31668 6666 31720 6672
rect 31772 6718 31892 6746
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 31680 6322 31708 6666
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31772 5914 31800 6718
rect 31852 6656 31904 6662
rect 31852 6598 31904 6604
rect 31864 6458 31892 6598
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31772 5030 31800 5850
rect 31852 5364 31904 5370
rect 31852 5306 31904 5312
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 31680 4622 31708 4966
rect 31772 4826 31800 4966
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31864 4486 31892 5306
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31404 3998 31524 4026
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31116 3460 31168 3466
rect 31116 3402 31168 3408
rect 31404 2990 31432 3998
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31496 3466 31524 3878
rect 31484 3460 31536 3466
rect 31484 3402 31536 3408
rect 31956 3058 31984 5170
rect 32048 4826 32076 7754
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 32140 7206 32168 7686
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32140 5302 32168 7142
rect 32232 6730 32260 9046
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32324 7546 32352 8910
rect 32312 7540 32364 7546
rect 32312 7482 32364 7488
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32220 6724 32272 6730
rect 32220 6666 32272 6672
rect 32416 6390 32444 7142
rect 32404 6384 32456 6390
rect 32404 6326 32456 6332
rect 32128 5296 32180 5302
rect 32128 5238 32180 5244
rect 32416 5250 32444 6326
rect 32508 6186 32536 9318
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32772 8832 32824 8838
rect 32772 8774 32824 8780
rect 32784 7478 32812 8774
rect 32864 8288 32916 8294
rect 32864 8230 32916 8236
rect 32772 7472 32824 7478
rect 32772 7414 32824 7420
rect 32588 6384 32640 6390
rect 32588 6326 32640 6332
rect 32496 6180 32548 6186
rect 32496 6122 32548 6128
rect 32600 5778 32628 6326
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32496 5296 32548 5302
rect 32416 5244 32496 5250
rect 32416 5238 32548 5244
rect 32416 5222 32536 5238
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 32600 4826 32628 4966
rect 32036 4820 32088 4826
rect 32036 4762 32088 4768
rect 32588 4820 32640 4826
rect 32588 4762 32640 4768
rect 32220 4752 32272 4758
rect 32220 4694 32272 4700
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 32140 3534 32168 4014
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32140 3058 32168 3470
rect 32232 3126 32260 4694
rect 32496 4548 32548 4554
rect 32496 4490 32548 4496
rect 32312 4480 32364 4486
rect 32312 4422 32364 4428
rect 32324 4146 32352 4422
rect 32508 4146 32536 4490
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32324 3534 32352 4082
rect 32508 3738 32536 4082
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 32876 3602 32904 8230
rect 32968 6458 32996 8910
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33048 8084 33100 8090
rect 33048 8026 33100 8032
rect 32956 6452 33008 6458
rect 32956 6394 33008 6400
rect 33060 5658 33088 8026
rect 33140 8016 33192 8022
rect 33140 7958 33192 7964
rect 32968 5642 33088 5658
rect 32956 5636 33088 5642
rect 33008 5630 33088 5636
rect 32956 5578 33008 5584
rect 33060 5370 33088 5630
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 33060 4554 33088 5306
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32876 3126 32904 3334
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 32864 3120 32916 3126
rect 32864 3062 32916 3068
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 31392 2984 31444 2990
rect 31392 2926 31444 2932
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 32036 2644 32088 2650
rect 32036 2586 32088 2592
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 30932 2100 30984 2106
rect 30932 2042 30984 2048
rect 31312 800 31340 2246
rect 32048 800 32076 2586
rect 32784 800 32812 2790
rect 33152 2446 33180 7958
rect 33244 7818 33272 8434
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33232 7812 33284 7818
rect 33232 7754 33284 7760
rect 33244 6390 33272 7754
rect 33232 6384 33284 6390
rect 33232 6326 33284 6332
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 33244 5098 33272 5646
rect 33336 5370 33364 7822
rect 33428 6458 33456 8434
rect 33416 6452 33468 6458
rect 33416 6394 33468 6400
rect 33428 6254 33456 6394
rect 33416 6248 33468 6254
rect 33416 6190 33468 6196
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 33232 5092 33284 5098
rect 33232 5034 33284 5040
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33428 4486 33456 4558
rect 33232 4480 33284 4486
rect 33232 4422 33284 4428
rect 33416 4480 33468 4486
rect 33416 4422 33468 4428
rect 33244 4282 33272 4422
rect 33232 4276 33284 4282
rect 33232 4218 33284 4224
rect 33324 4140 33376 4146
rect 33324 4082 33376 4088
rect 33336 3534 33364 4082
rect 33520 4026 33548 9318
rect 33612 7410 33640 9522
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33784 8628 33836 8634
rect 33784 8570 33836 8576
rect 33692 7744 33744 7750
rect 33692 7686 33744 7692
rect 33600 7404 33652 7410
rect 33600 7346 33652 7352
rect 33600 6656 33652 6662
rect 33600 6598 33652 6604
rect 33612 5642 33640 6598
rect 33600 5636 33652 5642
rect 33600 5578 33652 5584
rect 33600 4616 33652 4622
rect 33600 4558 33652 4564
rect 33428 4010 33548 4026
rect 33416 4004 33548 4010
rect 33468 3998 33548 4004
rect 33416 3946 33468 3952
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 33508 3460 33560 3466
rect 33508 3402 33560 3408
rect 33520 3194 33548 3402
rect 33508 3188 33560 3194
rect 33508 3130 33560 3136
rect 33612 3058 33640 4558
rect 33704 3058 33732 7686
rect 33796 6118 33824 8570
rect 33784 6112 33836 6118
rect 33784 6054 33836 6060
rect 33796 5914 33824 6054
rect 33888 5914 33916 8910
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 34520 8356 34572 8362
rect 34520 8298 34572 8304
rect 33968 7336 34020 7342
rect 33968 7278 34020 7284
rect 33980 6730 34008 7278
rect 33968 6724 34020 6730
rect 33968 6666 34020 6672
rect 33784 5908 33836 5914
rect 33784 5850 33836 5856
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 33968 5228 34020 5234
rect 33968 5170 34020 5176
rect 33980 4690 34008 5170
rect 33968 4684 34020 4690
rect 33968 4626 34020 4632
rect 33968 3732 34020 3738
rect 34072 3720 34100 8298
rect 34244 6452 34296 6458
rect 34244 6394 34296 6400
rect 34152 6384 34204 6390
rect 34152 6326 34204 6332
rect 34164 3738 34192 6326
rect 34256 4486 34284 6394
rect 34336 6180 34388 6186
rect 34336 6122 34388 6128
rect 34348 5098 34376 6122
rect 34428 6112 34480 6118
rect 34428 6054 34480 6060
rect 34440 5914 34468 6054
rect 34428 5908 34480 5914
rect 34428 5850 34480 5856
rect 34336 5092 34388 5098
rect 34336 5034 34388 5040
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34244 4480 34296 4486
rect 34244 4422 34296 4428
rect 34020 3692 34100 3720
rect 34152 3732 34204 3738
rect 33968 3674 34020 3680
rect 34152 3674 34204 3680
rect 34336 3664 34388 3670
rect 34336 3606 34388 3612
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 34348 2854 34376 3606
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 33508 2576 33560 2582
rect 33508 2518 33560 2524
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 33520 800 33548 2518
rect 34440 2514 34468 4966
rect 34532 4146 34560 8298
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34716 7478 34744 7686
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34808 7410 34836 7822
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34716 6254 34744 6734
rect 34808 6730 34836 7346
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34796 6724 34848 6730
rect 34796 6666 34848 6672
rect 34808 6322 34836 6666
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34624 4826 34652 5850
rect 34716 5166 34744 6190
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 34704 5160 34756 5166
rect 34704 5102 34756 5108
rect 34612 4820 34664 4826
rect 34612 4762 34664 4768
rect 34612 4276 34664 4282
rect 34612 4218 34664 4224
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 34624 3534 34652 4218
rect 34716 3942 34744 5102
rect 34808 4706 34836 5510
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35360 4826 35388 8434
rect 36084 7948 36136 7954
rect 36084 7890 36136 7896
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35440 7744 35492 7750
rect 35440 7686 35492 7692
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 35452 7206 35480 7686
rect 35440 7200 35492 7206
rect 35440 7142 35492 7148
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 34808 4678 34928 4706
rect 34900 4554 34928 4678
rect 34796 4548 34848 4554
rect 34796 4490 34848 4496
rect 34888 4548 34940 4554
rect 34888 4490 34940 4496
rect 34808 3942 34836 4490
rect 35452 4214 35480 7142
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35440 4208 35492 4214
rect 35440 4150 35492 4156
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 34716 3602 34744 3878
rect 34704 3596 34756 3602
rect 34704 3538 34756 3544
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 34624 3194 34652 3470
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 34808 3126 34836 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35452 3738 35480 3878
rect 35440 3732 35492 3738
rect 35440 3674 35492 3680
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34980 2576 35032 2582
rect 34980 2518 35032 2524
rect 34428 2508 34480 2514
rect 34428 2450 34480 2456
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 34256 800 34284 2246
rect 34992 800 35020 2518
rect 35544 2378 35572 5510
rect 35636 3466 35664 7686
rect 35728 4842 35756 7822
rect 36096 7478 36124 7890
rect 36452 7880 36504 7886
rect 36452 7822 36504 7828
rect 36636 7880 36688 7886
rect 36636 7822 36688 7828
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 36084 7472 36136 7478
rect 36084 7414 36136 7420
rect 36176 7404 36228 7410
rect 36176 7346 36228 7352
rect 35808 7200 35860 7206
rect 35808 7142 35860 7148
rect 35820 6390 35848 7142
rect 35900 6656 35952 6662
rect 35900 6598 35952 6604
rect 35808 6384 35860 6390
rect 35808 6326 35860 6332
rect 35728 4826 35848 4842
rect 35728 4820 35860 4826
rect 35728 4814 35808 4820
rect 35808 4762 35860 4768
rect 35624 3460 35676 3466
rect 35624 3402 35676 3408
rect 35912 3126 35940 6598
rect 36188 6458 36216 7346
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 36084 5704 36136 5710
rect 36084 5646 36136 5652
rect 35992 5568 36044 5574
rect 35992 5510 36044 5516
rect 35900 3120 35952 3126
rect 35900 3062 35952 3068
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 35532 2372 35584 2378
rect 35532 2314 35584 2320
rect 35728 800 35756 2858
rect 36004 2514 36032 5510
rect 36096 4690 36124 5646
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 36188 4554 36216 6394
rect 36280 5302 36308 7686
rect 36360 6112 36412 6118
rect 36360 6054 36412 6060
rect 36268 5296 36320 5302
rect 36268 5238 36320 5244
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 36176 4548 36228 4554
rect 36176 4490 36228 4496
rect 36096 3738 36124 4490
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 36096 3466 36124 3674
rect 36084 3460 36136 3466
rect 36084 3402 36136 3408
rect 35992 2508 36044 2514
rect 35992 2450 36044 2456
rect 36372 2446 36400 6054
rect 36464 5914 36492 7822
rect 36452 5908 36504 5914
rect 36452 5850 36504 5856
rect 36544 5636 36596 5642
rect 36544 5578 36596 5584
rect 36556 5370 36584 5578
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36544 5228 36596 5234
rect 36544 5170 36596 5176
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36464 4826 36492 4966
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36556 4622 36584 5170
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36452 3664 36504 3670
rect 36452 3606 36504 3612
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36464 800 36492 3606
rect 36648 3194 36676 7822
rect 37648 7744 37700 7750
rect 37648 7686 37700 7692
rect 37832 7744 37884 7750
rect 37832 7686 37884 7692
rect 36820 7404 36872 7410
rect 36820 7346 36872 7352
rect 36912 7404 36964 7410
rect 36912 7346 36964 7352
rect 36728 7268 36780 7274
rect 36728 7210 36780 7216
rect 36740 4146 36768 7210
rect 36832 6798 36860 7346
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 36820 6248 36872 6254
rect 36820 6190 36872 6196
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 36728 3392 36780 3398
rect 36728 3334 36780 3340
rect 36636 3188 36688 3194
rect 36636 3130 36688 3136
rect 36740 3058 36768 3334
rect 36832 3126 36860 6190
rect 36924 3738 36952 7346
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37188 6792 37240 6798
rect 37188 6734 37240 6740
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 36820 3120 36872 3126
rect 36820 3062 36872 3068
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 37108 2514 37136 5510
rect 37200 4078 37228 6734
rect 37292 4146 37320 7142
rect 37372 6656 37424 6662
rect 37372 6598 37424 6604
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37188 4072 37240 4078
rect 37188 4014 37240 4020
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 37096 2508 37148 2514
rect 37096 2450 37148 2456
rect 37200 800 37228 3878
rect 37384 3534 37412 6598
rect 37464 6112 37516 6118
rect 37464 6054 37516 6060
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37476 3058 37504 6054
rect 37660 4622 37688 7686
rect 37844 5710 37872 7686
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 38028 4826 38056 7822
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38120 5370 38148 7346
rect 39396 5568 39448 5574
rect 39396 5510 39448 5516
rect 38108 5364 38160 5370
rect 38108 5306 38160 5312
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 37648 4616 37700 4622
rect 37648 4558 37700 4564
rect 37924 4480 37976 4486
rect 37924 4422 37976 4428
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37936 800 37964 4422
rect 38660 4004 38712 4010
rect 38660 3946 38712 3952
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 2038 38056 2246
rect 38016 2032 38068 2038
rect 38016 1974 38068 1980
rect 38672 800 38700 3946
rect 39408 800 39436 5510
rect 39764 2372 39816 2378
rect 39764 2314 39816 2320
rect 39776 800 39804 2314
rect 23952 734 24164 762
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3974 9016 4030 9072
rect 3238 8472 3294 8528
rect 3606 8336 3662 8392
rect 202 3304 258 3360
rect 1674 6452 1730 6488
rect 1674 6432 1676 6452
rect 1676 6432 1728 6452
rect 1728 6432 1730 6452
rect 1858 5072 1914 5128
rect 2318 7656 2374 7712
rect 1674 3032 1730 3088
rect 2502 5480 2558 5536
rect 3238 7404 3294 7440
rect 3238 7384 3240 7404
rect 3240 7384 3292 7404
rect 3292 7384 3294 7404
rect 3146 5344 3202 5400
rect 2870 4140 2926 4176
rect 2870 4120 2872 4140
rect 2872 4120 2924 4140
rect 2924 4120 2926 4140
rect 3238 4664 3294 4720
rect 3422 5208 3478 5264
rect 3330 4392 3386 4448
rect 3330 4120 3386 4176
rect 3146 3188 3202 3224
rect 3146 3168 3148 3188
rect 3148 3168 3200 3188
rect 3200 3168 3202 3188
rect 3146 2896 3202 2952
rect 3422 3576 3478 3632
rect 3698 7540 3754 7576
rect 3698 7520 3700 7540
rect 3700 7520 3752 7540
rect 3752 7520 3754 7540
rect 3698 6332 3700 6352
rect 3700 6332 3752 6352
rect 3752 6332 3754 6352
rect 3698 6296 3754 6332
rect 3698 6160 3754 6216
rect 3698 5616 3754 5672
rect 4158 8744 4214 8800
rect 4066 8628 4122 8664
rect 4066 8608 4068 8628
rect 4068 8608 4120 8628
rect 4120 8608 4122 8628
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5078 8064 5134 8120
rect 4526 7828 4528 7848
rect 4528 7828 4580 7848
rect 4580 7828 4582 7848
rect 4526 7792 4582 7828
rect 3790 4548 3846 4584
rect 3790 4528 3792 4548
rect 3792 4528 3844 4548
rect 3844 4528 3846 4548
rect 3606 3984 3662 4040
rect 3790 3440 3846 3496
rect 4434 7248 4490 7304
rect 4894 7148 4896 7168
rect 4896 7148 4948 7168
rect 4948 7148 4950 7168
rect 4894 7112 4950 7148
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 5354 7656 5410 7712
rect 5354 6840 5410 6896
rect 5078 6024 5134 6080
rect 4986 5752 5042 5808
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4894 5208 4950 5264
rect 4894 3848 4950 3904
rect 5998 8084 6054 8120
rect 5998 8064 6000 8084
rect 6000 8064 6052 8084
rect 6052 8064 6054 8084
rect 5538 3712 5594 3768
rect 5906 3848 5962 3904
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6182 3712 6238 3768
rect 7470 9016 7526 9072
rect 6918 8472 6974 8528
rect 6366 4528 6422 4584
rect 7010 8336 7066 8392
rect 6642 6432 6698 6488
rect 6918 6432 6974 6488
rect 7010 5480 7066 5536
rect 7470 5480 7526 5536
rect 7194 3068 7196 3088
rect 7196 3068 7248 3088
rect 7248 3068 7250 3088
rect 7194 3032 7250 3068
rect 9310 8608 9366 8664
rect 7838 7520 7894 7576
rect 8298 7112 8354 7168
rect 8390 6196 8392 6216
rect 8392 6196 8444 6216
rect 8444 6196 8446 6216
rect 8390 6160 8446 6196
rect 8298 6024 8354 6080
rect 8298 3848 8354 3904
rect 7470 3032 7526 3088
rect 8390 3576 8446 3632
rect 8666 5788 8668 5808
rect 8668 5788 8720 5808
rect 8720 5788 8722 5808
rect 8666 5752 8722 5788
rect 8574 3188 8630 3224
rect 8574 3168 8576 3188
rect 8576 3168 8628 3188
rect 8628 3168 8630 3188
rect 8942 6432 8998 6488
rect 9494 6840 9550 6896
rect 10046 8916 10048 8936
rect 10048 8916 10100 8936
rect 10100 8916 10102 8936
rect 10046 8880 10102 8916
rect 10414 8744 10470 8800
rect 9678 7792 9734 7848
rect 9770 7248 9826 7304
rect 9678 6316 9734 6352
rect 9678 6296 9680 6316
rect 9680 6296 9732 6316
rect 9732 6296 9734 6316
rect 9770 4936 9826 4992
rect 10322 6160 10378 6216
rect 10230 5480 10286 5536
rect 9862 4664 9918 4720
rect 8942 4120 8998 4176
rect 9678 4156 9680 4176
rect 9680 4156 9732 4176
rect 9732 4156 9734 4176
rect 9678 4120 9734 4156
rect 9126 3052 9182 3088
rect 9126 3032 9128 3052
rect 9128 3032 9180 3052
rect 9180 3032 9182 3052
rect 9310 2896 9366 2952
rect 10414 4800 10470 4856
rect 10782 9596 10784 9616
rect 10784 9596 10836 9616
rect 10836 9596 10838 9616
rect 10782 9560 10838 9596
rect 10598 3576 10654 3632
rect 10874 5616 10930 5672
rect 10966 5480 11022 5536
rect 10966 4800 11022 4856
rect 11058 4256 11114 4312
rect 11334 5344 11390 5400
rect 12530 8744 12586 8800
rect 11518 7384 11574 7440
rect 11426 5072 11482 5128
rect 11886 6296 11942 6352
rect 11518 4256 11574 4312
rect 11978 4392 12034 4448
rect 11978 4276 12034 4312
rect 11978 4256 11980 4276
rect 11980 4256 12032 4276
rect 12032 4256 12034 4276
rect 11978 3848 12034 3904
rect 12622 6316 12678 6352
rect 12622 6296 12624 6316
rect 12624 6296 12676 6316
rect 12676 6296 12678 6316
rect 13266 9560 13322 9616
rect 14002 13268 14004 13288
rect 14004 13268 14056 13288
rect 14056 13268 14058 13288
rect 14002 13232 14058 13268
rect 12622 5480 12678 5536
rect 12254 3732 12310 3768
rect 12254 3712 12256 3732
rect 12256 3712 12308 3732
rect 12308 3712 12310 3732
rect 12346 3576 12402 3632
rect 12714 3984 12770 4040
rect 13450 9016 13506 9072
rect 13634 7248 13690 7304
rect 13174 3460 13230 3496
rect 13174 3440 13176 3460
rect 13176 3440 13228 3460
rect 13228 3440 13230 3460
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 14186 4140 14242 4176
rect 14186 4120 14188 4140
rect 14188 4120 14240 4140
rect 14240 4120 14242 4140
rect 14278 3576 14334 3632
rect 15382 12824 15438 12880
rect 15106 11056 15162 11112
rect 14646 3984 14702 4040
rect 15382 8880 15438 8936
rect 15014 7248 15070 7304
rect 15382 6840 15438 6896
rect 15566 7248 15622 7304
rect 14830 3576 14886 3632
rect 15474 4972 15476 4992
rect 15476 4972 15528 4992
rect 15528 4972 15530 4992
rect 15474 4936 15530 4972
rect 16854 15816 16910 15872
rect 16670 11192 16726 11248
rect 16302 6160 16358 6216
rect 16946 10920 17002 10976
rect 16946 9424 17002 9480
rect 16854 9152 16910 9208
rect 16670 4120 16726 4176
rect 16762 3712 16818 3768
rect 17038 3884 17040 3904
rect 17040 3884 17092 3904
rect 17092 3884 17094 3904
rect 17038 3848 17094 3884
rect 19982 28328 20038 28384
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 17774 17448 17830 17504
rect 17682 15816 17738 15872
rect 17222 9324 17224 9344
rect 17224 9324 17276 9344
rect 17276 9324 17278 9344
rect 17222 9288 17278 9324
rect 17498 9560 17554 9616
rect 17590 6704 17646 6760
rect 17866 10920 17922 10976
rect 18694 13776 18750 13832
rect 18510 11192 18566 11248
rect 18326 8744 18382 8800
rect 18602 9172 18658 9208
rect 18602 9152 18604 9172
rect 18604 9152 18656 9172
rect 18656 9152 18658 9172
rect 18418 8608 18474 8664
rect 18234 3596 18290 3632
rect 18234 3576 18236 3596
rect 18236 3576 18288 3596
rect 18288 3576 18290 3596
rect 19982 27276 19984 27296
rect 19984 27276 20036 27296
rect 20036 27276 20038 27296
rect 19982 27240 20038 27276
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19890 24248 19946 24304
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19890 23060 19892 23080
rect 19892 23060 19944 23080
rect 19944 23060 19946 23080
rect 19890 23024 19946 23060
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20074 22480 20130 22536
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20350 22208 20406 22264
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20074 19760 20130 19816
rect 19982 19488 20038 19544
rect 19430 18808 19486 18864
rect 19798 18692 19854 18728
rect 19798 18672 19800 18692
rect 19800 18672 19852 18692
rect 19852 18672 19854 18692
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19522 18128 19578 18184
rect 19614 17720 19670 17776
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19522 16632 19578 16688
rect 19522 16532 19524 16552
rect 19524 16532 19576 16552
rect 19576 16532 19578 16552
rect 19522 16496 19578 16532
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19706 15952 19762 16008
rect 19614 15680 19670 15736
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19522 14900 19524 14920
rect 19524 14900 19576 14920
rect 19576 14900 19578 14920
rect 19522 14864 19578 14900
rect 19890 14592 19946 14648
rect 19338 13912 19394 13968
rect 19154 13640 19210 13696
rect 18878 9036 18934 9072
rect 18878 9016 18880 9036
rect 18880 9016 18932 9036
rect 18932 9016 18934 9036
rect 19062 9460 19064 9480
rect 19064 9460 19116 9480
rect 19116 9460 19118 9480
rect 19062 9424 19118 9460
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 21822 28364 21824 28384
rect 21824 28364 21876 28384
rect 21876 28364 21878 28384
rect 21822 28328 21878 28364
rect 20718 19932 20720 19952
rect 20720 19932 20772 19952
rect 20772 19932 20774 19952
rect 20718 19896 20774 19932
rect 20810 19760 20866 19816
rect 20718 18672 20774 18728
rect 21178 19488 21234 19544
rect 20994 18708 20996 18728
rect 20996 18708 21048 18728
rect 21048 18708 21050 18728
rect 20994 18672 21050 18708
rect 20902 18536 20958 18592
rect 20902 18284 20958 18320
rect 20902 18264 20904 18284
rect 20904 18264 20956 18284
rect 20956 18264 20958 18284
rect 20350 13776 20406 13832
rect 19522 13368 19578 13424
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19246 10668 19302 10704
rect 19246 10648 19248 10668
rect 19248 10648 19300 10668
rect 19300 10648 19302 10668
rect 20350 13368 20406 13424
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19982 9288 20038 9344
rect 19522 9152 19578 9208
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19430 8628 19486 8664
rect 19430 8608 19432 8628
rect 19432 8608 19484 8628
rect 19484 8608 19486 8628
rect 19982 8472 20038 8528
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20258 10104 20314 10160
rect 20258 8608 20314 8664
rect 20534 14728 20590 14784
rect 21086 18264 21142 18320
rect 20994 15408 21050 15464
rect 21086 14864 21142 14920
rect 20534 13912 20590 13968
rect 20442 8336 20498 8392
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19890 6316 19946 6352
rect 19890 6296 19892 6316
rect 19892 6296 19944 6316
rect 19944 6296 19946 6316
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19154 3984 19210 4040
rect 19338 3576 19394 3632
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19614 4156 19616 4176
rect 19616 4156 19668 4176
rect 19668 4156 19670 4176
rect 19614 4120 19670 4156
rect 19522 3848 19578 3904
rect 19430 3440 19486 3496
rect 19798 3712 19854 3768
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19430 2896 19486 2952
rect 19798 2760 19854 2816
rect 20442 7384 20498 7440
rect 20626 11736 20682 11792
rect 20626 11464 20682 11520
rect 21086 14728 21142 14784
rect 20994 13776 21050 13832
rect 20994 13524 21050 13560
rect 20994 13504 20996 13524
rect 20996 13504 21048 13524
rect 21048 13504 21050 13524
rect 21454 19796 21456 19816
rect 21456 19796 21508 19816
rect 21508 19796 21510 19816
rect 21454 19760 21510 19796
rect 21638 20596 21694 20632
rect 21638 20576 21640 20596
rect 21640 20576 21692 20596
rect 21692 20576 21694 20596
rect 21638 18808 21694 18864
rect 21822 18536 21878 18592
rect 21362 16224 21418 16280
rect 21086 10920 21142 10976
rect 20810 8608 20866 8664
rect 20994 8744 21050 8800
rect 20534 6160 20590 6216
rect 20350 3984 20406 4040
rect 20258 3576 20314 3632
rect 19522 2488 19578 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20534 2896 20590 2952
rect 20994 6568 21050 6624
rect 20994 6316 21050 6352
rect 20994 6296 20996 6316
rect 20996 6296 21048 6316
rect 21048 6296 21050 6316
rect 20718 4140 20774 4176
rect 20718 4120 20720 4140
rect 20720 4120 20772 4140
rect 20772 4120 20774 4140
rect 20810 3576 20866 3632
rect 20994 3984 21050 4040
rect 21546 16360 21602 16416
rect 21730 16904 21786 16960
rect 21730 16768 21786 16824
rect 21546 15952 21602 16008
rect 21546 15544 21602 15600
rect 21546 14592 21602 14648
rect 23478 24248 23534 24304
rect 22926 23316 22982 23352
rect 22926 23296 22928 23316
rect 22928 23296 22980 23316
rect 22980 23296 22982 23316
rect 22650 21392 22706 21448
rect 22374 19896 22430 19952
rect 22466 18708 22468 18728
rect 22468 18708 22520 18728
rect 22520 18708 22522 18728
rect 22466 18672 22522 18708
rect 21914 15952 21970 16008
rect 22098 15952 22154 16008
rect 21730 13232 21786 13288
rect 21454 9968 21510 10024
rect 21730 10920 21786 10976
rect 22190 14592 22246 14648
rect 22098 14456 22154 14512
rect 22006 14220 22008 14240
rect 22008 14220 22060 14240
rect 22060 14220 22062 14240
rect 22006 14184 22062 14220
rect 22190 12688 22246 12744
rect 22466 14320 22522 14376
rect 22466 12552 22522 12608
rect 21822 9560 21878 9616
rect 21822 8880 21878 8936
rect 22374 9560 22430 9616
rect 22098 9324 22100 9344
rect 22100 9324 22152 9344
rect 22152 9324 22154 9344
rect 22098 9288 22154 9324
rect 22006 9016 22062 9072
rect 22006 8336 22062 8392
rect 22650 15680 22706 15736
rect 23386 18028 23388 18048
rect 23388 18028 23440 18048
rect 23440 18028 23442 18048
rect 23386 17992 23442 18028
rect 23110 14456 23166 14512
rect 22742 12552 22798 12608
rect 22834 11736 22890 11792
rect 22650 9560 22706 9616
rect 22650 9016 22706 9072
rect 23110 11600 23166 11656
rect 23202 11192 23258 11248
rect 22926 10240 22982 10296
rect 22926 10104 22982 10160
rect 23018 8372 23020 8392
rect 23020 8372 23072 8392
rect 23072 8372 23074 8392
rect 23018 8336 23074 8372
rect 22926 7656 22982 7712
rect 22374 6316 22430 6352
rect 22374 6296 22376 6316
rect 22376 6296 22428 6316
rect 22428 6296 22430 6316
rect 23478 14184 23534 14240
rect 23386 10240 23442 10296
rect 23294 8336 23350 8392
rect 23294 7248 23350 7304
rect 24030 23432 24086 23488
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 25226 23432 25282 23488
rect 25318 22072 25374 22128
rect 25502 23296 25558 23352
rect 24950 19216 25006 19272
rect 25042 16904 25098 16960
rect 24674 16496 24730 16552
rect 24214 15020 24270 15056
rect 24214 15000 24216 15020
rect 24216 15000 24268 15020
rect 24268 15000 24270 15020
rect 24122 14900 24124 14920
rect 24124 14900 24176 14920
rect 24176 14900 24178 14920
rect 24122 14864 24178 14900
rect 24030 13640 24086 13696
rect 24950 15816 25006 15872
rect 24398 14764 24400 14784
rect 24400 14764 24452 14784
rect 24452 14764 24454 14784
rect 24398 14728 24454 14764
rect 24122 12708 24178 12744
rect 24122 12688 24124 12708
rect 24124 12688 24176 12708
rect 24176 12688 24178 12708
rect 23570 10920 23626 10976
rect 23938 10648 23994 10704
rect 23478 6024 23534 6080
rect 23386 5908 23442 5944
rect 23386 5888 23388 5908
rect 23388 5888 23440 5908
rect 23440 5888 23442 5908
rect 23294 3848 23350 3904
rect 23478 3712 23534 3768
rect 24030 9560 24086 9616
rect 24950 15136 25006 15192
rect 24858 14728 24914 14784
rect 24674 9580 24730 9616
rect 24674 9560 24676 9580
rect 24676 9560 24728 9580
rect 24728 9560 24730 9580
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 25318 14864 25374 14920
rect 25686 15136 25742 15192
rect 25686 13640 25742 13696
rect 25502 11056 25558 11112
rect 25042 8628 25098 8664
rect 25042 8608 25044 8628
rect 25044 8608 25096 8628
rect 25096 8608 25098 8628
rect 24306 6296 24362 6352
rect 25962 15000 26018 15056
rect 26146 15680 26202 15736
rect 26422 18128 26478 18184
rect 26330 11328 26386 11384
rect 25962 11192 26018 11248
rect 26514 11600 26570 11656
rect 26054 10920 26110 10976
rect 25686 9596 25688 9616
rect 25688 9596 25740 9616
rect 25740 9596 25742 9616
rect 25686 9560 25742 9596
rect 25134 6060 25136 6080
rect 25136 6060 25188 6080
rect 25188 6060 25190 6080
rect 25134 6024 25190 6060
rect 25778 5752 25834 5808
rect 25686 3848 25742 3904
rect 27526 21664 27582 21720
rect 27066 15408 27122 15464
rect 26790 14320 26846 14376
rect 26698 10920 26754 10976
rect 26514 9424 26570 9480
rect 26882 10784 26938 10840
rect 28262 21140 28318 21176
rect 28262 21120 28264 21140
rect 28264 21120 28316 21140
rect 28316 21120 28318 21140
rect 29182 21548 29238 21584
rect 29182 21528 29184 21548
rect 29184 21528 29236 21548
rect 29236 21528 29238 21548
rect 28814 21392 28870 21448
rect 28998 21392 29054 21448
rect 28814 21120 28870 21176
rect 30010 23060 30012 23080
rect 30012 23060 30064 23080
rect 30064 23060 30066 23080
rect 30010 23024 30066 23060
rect 29918 21936 29974 21992
rect 31206 23044 31262 23080
rect 31206 23024 31208 23044
rect 31208 23024 31260 23044
rect 31260 23024 31262 23044
rect 27802 15544 27858 15600
rect 27066 8900 27122 8936
rect 27066 8880 27068 8900
rect 27068 8880 27120 8900
rect 27120 8880 27122 8900
rect 27526 11056 27582 11112
rect 27802 10920 27858 10976
rect 27986 12280 28042 12336
rect 27710 9424 27766 9480
rect 27618 9152 27674 9208
rect 27526 9016 27582 9072
rect 26882 5636 26938 5672
rect 26882 5616 26884 5636
rect 26884 5616 26936 5636
rect 26936 5616 26938 5636
rect 27434 7656 27490 7712
rect 27434 5772 27490 5808
rect 27434 5752 27436 5772
rect 27436 5752 27488 5772
rect 27488 5752 27490 5772
rect 27894 9288 27950 9344
rect 28630 19236 28686 19272
rect 28630 19216 28632 19236
rect 28632 19216 28684 19236
rect 28684 19216 28686 19236
rect 28170 12280 28226 12336
rect 28170 8608 28226 8664
rect 30746 21392 30802 21448
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35622 21936 35678 21992
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 28722 10648 28778 10704
rect 28538 8880 28594 8936
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 28262 7384 28318 7440
rect 27986 7248 28042 7304
rect 27986 5888 28042 5944
rect 28078 5616 28134 5672
rect 28170 4140 28226 4176
rect 28170 4120 28172 4140
rect 28172 4120 28224 4140
rect 28224 4120 28226 4140
rect 31482 11192 31538 11248
rect 29550 9832 29606 9888
rect 29090 8744 29146 8800
rect 28814 4140 28870 4176
rect 28814 4120 28816 4140
rect 28816 4120 28868 4140
rect 28868 4120 28870 4140
rect 29918 6704 29974 6760
rect 30746 9832 30802 9888
rect 30562 9424 30618 9480
rect 30654 9016 30710 9072
rect 28722 2760 28778 2816
rect 31298 6840 31354 6896
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 31482 6840 31538 6896
rect 31758 6840 31814 6896
rect 31942 7520 31998 7576
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19977 28386 20043 28389
rect 21817 28386 21883 28389
rect 19977 28384 21883 28386
rect 19977 28328 19982 28384
rect 20038 28328 21822 28384
rect 21878 28328 21883 28384
rect 19977 28326 21883 28328
rect 19977 28323 20043 28326
rect 21817 28323 21883 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19977 27298 20043 27301
rect 20294 27298 20300 27300
rect 19977 27296 20300 27298
rect 19977 27240 19982 27296
rect 20038 27240 20300 27296
rect 19977 27238 20300 27240
rect 19977 27235 20043 27238
rect 20294 27236 20300 27238
rect 20364 27236 20370 27300
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 19885 24306 19951 24309
rect 23473 24306 23539 24309
rect 19885 24304 23539 24306
rect 19885 24248 19890 24304
rect 19946 24248 23478 24304
rect 23534 24248 23539 24304
rect 19885 24246 23539 24248
rect 19885 24243 19951 24246
rect 23473 24243 23539 24246
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 24025 23490 24091 23493
rect 25221 23490 25287 23493
rect 24025 23488 25287 23490
rect 24025 23432 24030 23488
rect 24086 23432 25226 23488
rect 25282 23432 25287 23488
rect 24025 23430 25287 23432
rect 24025 23427 24091 23430
rect 25221 23427 25287 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 22921 23354 22987 23357
rect 25497 23354 25563 23357
rect 22921 23352 25563 23354
rect 22921 23296 22926 23352
rect 22982 23296 25502 23352
rect 25558 23296 25563 23352
rect 22921 23294 25563 23296
rect 22921 23291 22987 23294
rect 25497 23291 25563 23294
rect 19885 23082 19951 23085
rect 30005 23082 30071 23085
rect 31201 23082 31267 23085
rect 19885 23080 20178 23082
rect 19885 23024 19890 23080
rect 19946 23024 20178 23080
rect 19885 23022 20178 23024
rect 19885 23019 19951 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 20118 22541 20178 23022
rect 30005 23080 31267 23082
rect 30005 23024 30010 23080
rect 30066 23024 31206 23080
rect 31262 23024 31267 23080
rect 30005 23022 31267 23024
rect 30005 23019 30071 23022
rect 31201 23019 31267 23022
rect 20069 22536 20178 22541
rect 20069 22480 20074 22536
rect 20130 22480 20178 22536
rect 20069 22478 20178 22480
rect 20069 22475 20135 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 20345 22268 20411 22269
rect 20294 22266 20300 22268
rect 20254 22206 20300 22266
rect 20364 22264 20411 22268
rect 20406 22208 20411 22264
rect 20294 22204 20300 22206
rect 20364 22204 20411 22208
rect 20345 22203 20411 22204
rect 25313 22130 25379 22133
rect 25313 22128 29010 22130
rect 25313 22072 25318 22128
rect 25374 22072 29010 22128
rect 25313 22070 29010 22072
rect 25313 22067 25379 22070
rect 28950 21994 29010 22070
rect 29913 21994 29979 21997
rect 35617 21994 35683 21997
rect 28950 21992 35683 21994
rect 28950 21936 29918 21992
rect 29974 21936 35622 21992
rect 35678 21936 35683 21992
rect 28950 21934 35683 21936
rect 29913 21931 29979 21934
rect 35617 21931 35683 21934
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 27521 21722 27587 21725
rect 27521 21720 28872 21722
rect 27521 21664 27526 21720
rect 27582 21664 28872 21720
rect 27521 21662 28872 21664
rect 27521 21659 27587 21662
rect 28812 21586 28872 21662
rect 29177 21586 29243 21589
rect 28812 21584 29243 21586
rect 28812 21528 29182 21584
rect 29238 21528 29243 21584
rect 28812 21526 29243 21528
rect 29177 21523 29243 21526
rect 22645 21450 22711 21453
rect 28809 21450 28875 21453
rect 22645 21448 28875 21450
rect 22645 21392 22650 21448
rect 22706 21392 28814 21448
rect 28870 21392 28875 21448
rect 22645 21390 28875 21392
rect 22645 21387 22711 21390
rect 28809 21387 28875 21390
rect 28993 21450 29059 21453
rect 30741 21450 30807 21453
rect 28993 21448 30807 21450
rect 28993 21392 28998 21448
rect 29054 21392 30746 21448
rect 30802 21392 30807 21448
rect 28993 21390 30807 21392
rect 28993 21387 29059 21390
rect 30741 21387 30807 21390
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 28257 21178 28323 21181
rect 28809 21178 28875 21181
rect 28257 21176 28875 21178
rect 28257 21120 28262 21176
rect 28318 21120 28814 21176
rect 28870 21120 28875 21176
rect 28257 21118 28875 21120
rect 28257 21115 28323 21118
rect 28809 21115 28875 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 21633 20636 21699 20637
rect 21582 20634 21588 20636
rect 21542 20574 21588 20634
rect 21652 20632 21699 20636
rect 21694 20576 21699 20632
rect 21582 20572 21588 20574
rect 21652 20572 21699 20576
rect 21633 20571 21699 20572
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 20713 19954 20779 19957
rect 22369 19954 22435 19957
rect 20713 19952 22435 19954
rect 20713 19896 20718 19952
rect 20774 19896 22374 19952
rect 22430 19896 22435 19952
rect 20713 19894 22435 19896
rect 20713 19891 20779 19894
rect 22369 19891 22435 19894
rect 20069 19818 20135 19821
rect 20805 19818 20871 19821
rect 21449 19818 21515 19821
rect 20069 19816 21515 19818
rect 20069 19760 20074 19816
rect 20130 19760 20810 19816
rect 20866 19760 21454 19816
rect 21510 19760 21515 19816
rect 20069 19758 21515 19760
rect 20069 19755 20135 19758
rect 20805 19755 20871 19758
rect 21449 19755 21515 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 19977 19546 20043 19549
rect 21173 19546 21239 19549
rect 19977 19544 21239 19546
rect 19977 19488 19982 19544
rect 20038 19488 21178 19544
rect 21234 19488 21239 19544
rect 19977 19486 21239 19488
rect 19977 19483 20043 19486
rect 21173 19483 21239 19486
rect 24945 19274 25011 19277
rect 28625 19274 28691 19277
rect 24945 19272 28691 19274
rect 24945 19216 24950 19272
rect 25006 19216 28630 19272
rect 28686 19216 28691 19272
rect 24945 19214 28691 19216
rect 24945 19211 25011 19214
rect 28625 19211 28691 19214
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19425 18866 19491 18869
rect 21633 18866 21699 18869
rect 19425 18864 21699 18866
rect 19425 18808 19430 18864
rect 19486 18808 21638 18864
rect 21694 18808 21699 18864
rect 19425 18806 21699 18808
rect 19425 18803 19491 18806
rect 20670 18733 20730 18806
rect 21633 18803 21699 18806
rect 19793 18730 19859 18733
rect 20294 18730 20300 18732
rect 19793 18728 20300 18730
rect 19793 18672 19798 18728
rect 19854 18672 20300 18728
rect 19793 18670 20300 18672
rect 19793 18667 19859 18670
rect 20294 18668 20300 18670
rect 20364 18668 20370 18732
rect 20670 18728 20779 18733
rect 20670 18672 20718 18728
rect 20774 18672 20779 18728
rect 20670 18670 20779 18672
rect 20713 18667 20779 18670
rect 20989 18730 21055 18733
rect 22461 18730 22527 18733
rect 20989 18728 22527 18730
rect 20989 18672 20994 18728
rect 21050 18672 22466 18728
rect 22522 18672 22527 18728
rect 20989 18670 22527 18672
rect 20989 18667 21055 18670
rect 22461 18667 22527 18670
rect 20897 18594 20963 18597
rect 21030 18594 21036 18596
rect 20897 18592 21036 18594
rect 20897 18536 20902 18592
rect 20958 18536 21036 18592
rect 20897 18534 21036 18536
rect 20897 18531 20963 18534
rect 21030 18532 21036 18534
rect 21100 18532 21106 18596
rect 21817 18594 21883 18597
rect 21950 18594 21956 18596
rect 21817 18592 21956 18594
rect 21817 18536 21822 18592
rect 21878 18536 21956 18592
rect 21817 18534 21956 18536
rect 21817 18531 21883 18534
rect 21950 18532 21956 18534
rect 22020 18532 22026 18596
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 20897 18322 20963 18325
rect 21081 18322 21147 18325
rect 20897 18320 21147 18322
rect 20897 18264 20902 18320
rect 20958 18264 21086 18320
rect 21142 18264 21147 18320
rect 20897 18262 21147 18264
rect 20897 18259 20963 18262
rect 21081 18259 21147 18262
rect 19517 18186 19583 18189
rect 26417 18186 26483 18189
rect 19517 18184 26483 18186
rect 19517 18128 19522 18184
rect 19578 18128 26422 18184
rect 26478 18128 26483 18184
rect 19517 18126 26483 18128
rect 19517 18123 19583 18126
rect 26417 18123 26483 18126
rect 23238 17988 23244 18052
rect 23308 18050 23314 18052
rect 23381 18050 23447 18053
rect 23308 18048 23447 18050
rect 23308 17992 23386 18048
rect 23442 17992 23447 18048
rect 23308 17990 23447 17992
rect 23308 17988 23314 17990
rect 23381 17987 23447 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19609 17778 19675 17781
rect 19014 17776 19675 17778
rect 19014 17720 19614 17776
rect 19670 17720 19675 17776
rect 19014 17718 19675 17720
rect 17769 17506 17835 17509
rect 19014 17506 19074 17718
rect 19609 17715 19675 17718
rect 17769 17504 19074 17506
rect 17769 17448 17774 17504
rect 17830 17448 19074 17504
rect 17769 17446 19074 17448
rect 17769 17443 17835 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 21725 16962 21791 16965
rect 25037 16962 25103 16965
rect 21725 16960 25103 16962
rect 21725 16904 21730 16960
rect 21786 16904 25042 16960
rect 25098 16904 25103 16960
rect 21725 16902 25103 16904
rect 21725 16899 21791 16902
rect 25037 16899 25103 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 21030 16764 21036 16828
rect 21100 16826 21106 16828
rect 21725 16826 21791 16829
rect 21100 16824 21791 16826
rect 21100 16768 21730 16824
rect 21786 16768 21791 16824
rect 21100 16766 21791 16768
rect 21100 16764 21106 16766
rect 21725 16763 21791 16766
rect 19374 16628 19380 16692
rect 19444 16690 19450 16692
rect 19517 16690 19583 16693
rect 19444 16688 19583 16690
rect 19444 16632 19522 16688
rect 19578 16632 19583 16688
rect 19444 16630 19583 16632
rect 19444 16628 19450 16630
rect 19517 16627 19583 16630
rect 19517 16554 19583 16557
rect 20478 16554 20484 16556
rect 19517 16552 20484 16554
rect 19517 16496 19522 16552
rect 19578 16496 20484 16552
rect 19517 16494 20484 16496
rect 19517 16491 19583 16494
rect 20478 16492 20484 16494
rect 20548 16554 20554 16556
rect 24669 16554 24735 16557
rect 20548 16552 24735 16554
rect 20548 16496 24674 16552
rect 24730 16496 24735 16552
rect 20548 16494 24735 16496
rect 20548 16492 20554 16494
rect 24669 16491 24735 16494
rect 21541 16416 21607 16421
rect 21541 16360 21546 16416
rect 21602 16360 21607 16416
rect 21541 16355 21607 16360
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 21357 16282 21423 16285
rect 21544 16282 21604 16355
rect 21357 16280 21604 16282
rect 21357 16224 21362 16280
rect 21418 16224 21604 16280
rect 21357 16222 21604 16224
rect 21357 16219 21423 16222
rect 20110 16084 20116 16148
rect 20180 16146 20186 16148
rect 21582 16146 21588 16148
rect 20180 16086 21588 16146
rect 20180 16084 20186 16086
rect 21582 16084 21588 16086
rect 21652 16084 21658 16148
rect 19701 16010 19767 16013
rect 20846 16010 20852 16012
rect 19701 16008 20852 16010
rect 19701 15952 19706 16008
rect 19762 15952 20852 16008
rect 19701 15950 20852 15952
rect 19701 15947 19767 15950
rect 20846 15948 20852 15950
rect 20916 16010 20922 16012
rect 21541 16010 21607 16013
rect 20916 16008 21607 16010
rect 20916 15952 21546 16008
rect 21602 15952 21607 16008
rect 20916 15950 21607 15952
rect 20916 15948 20922 15950
rect 21541 15947 21607 15950
rect 21909 16010 21975 16013
rect 22093 16010 22159 16013
rect 21909 16008 22159 16010
rect 21909 15952 21914 16008
rect 21970 15952 22098 16008
rect 22154 15952 22159 16008
rect 21909 15950 22159 15952
rect 21909 15947 21975 15950
rect 22093 15947 22159 15950
rect 16849 15874 16915 15877
rect 17677 15874 17743 15877
rect 24945 15874 25011 15877
rect 16849 15872 25011 15874
rect 16849 15816 16854 15872
rect 16910 15816 17682 15872
rect 17738 15816 24950 15872
rect 25006 15816 25011 15872
rect 16849 15814 25011 15816
rect 16849 15811 16915 15814
rect 17677 15811 17743 15814
rect 24945 15811 25011 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19609 15738 19675 15741
rect 20110 15738 20116 15740
rect 19609 15736 20116 15738
rect 19609 15680 19614 15736
rect 19670 15680 20116 15736
rect 19609 15678 20116 15680
rect 19609 15675 19675 15678
rect 20110 15676 20116 15678
rect 20180 15676 20186 15740
rect 22645 15738 22711 15741
rect 26141 15738 26207 15741
rect 22645 15736 26207 15738
rect 22645 15680 22650 15736
rect 22706 15680 26146 15736
rect 26202 15680 26207 15736
rect 22645 15678 26207 15680
rect 22645 15675 22711 15678
rect 26141 15675 26207 15678
rect 21541 15602 21607 15605
rect 27797 15602 27863 15605
rect 21541 15600 27863 15602
rect 21541 15544 21546 15600
rect 21602 15544 27802 15600
rect 27858 15544 27863 15600
rect 21541 15542 27863 15544
rect 21541 15539 21607 15542
rect 27797 15539 27863 15542
rect 20989 15466 21055 15469
rect 27061 15466 27127 15469
rect 20989 15464 27127 15466
rect 20989 15408 20994 15464
rect 21050 15408 27066 15464
rect 27122 15408 27127 15464
rect 20989 15406 27127 15408
rect 20989 15403 21055 15406
rect 27061 15403 27127 15406
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 24945 15194 25011 15197
rect 25681 15194 25747 15197
rect 24945 15192 25747 15194
rect 24945 15136 24950 15192
rect 25006 15136 25686 15192
rect 25742 15136 25747 15192
rect 24945 15134 25747 15136
rect 24945 15131 25011 15134
rect 25681 15131 25747 15134
rect 24209 15058 24275 15061
rect 25957 15058 26023 15061
rect 24209 15056 26023 15058
rect 24209 15000 24214 15056
rect 24270 15000 25962 15056
rect 26018 15000 26023 15056
rect 24209 14998 26023 15000
rect 24209 14995 24275 14998
rect 25957 14995 26023 14998
rect 19190 14860 19196 14924
rect 19260 14922 19266 14924
rect 19517 14922 19583 14925
rect 21081 14922 21147 14925
rect 19260 14920 21147 14922
rect 19260 14864 19522 14920
rect 19578 14864 21086 14920
rect 21142 14864 21147 14920
rect 19260 14862 21147 14864
rect 19260 14860 19266 14862
rect 19517 14859 19583 14862
rect 21081 14859 21147 14862
rect 24117 14922 24183 14925
rect 25313 14922 25379 14925
rect 24117 14920 25379 14922
rect 24117 14864 24122 14920
rect 24178 14864 25318 14920
rect 25374 14864 25379 14920
rect 24117 14862 25379 14864
rect 24117 14859 24183 14862
rect 25313 14859 25379 14862
rect 20529 14786 20595 14789
rect 21081 14786 21147 14789
rect 20529 14784 21147 14786
rect 20529 14728 20534 14784
rect 20590 14728 21086 14784
rect 21142 14728 21147 14784
rect 20529 14726 21147 14728
rect 20529 14723 20595 14726
rect 21081 14723 21147 14726
rect 24393 14786 24459 14789
rect 24853 14786 24919 14789
rect 24393 14784 24919 14786
rect 24393 14728 24398 14784
rect 24454 14728 24858 14784
rect 24914 14728 24919 14784
rect 24393 14726 24919 14728
rect 24393 14723 24459 14726
rect 24853 14723 24919 14726
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19885 14650 19951 14653
rect 21541 14650 21607 14653
rect 19885 14648 21607 14650
rect 19885 14592 19890 14648
rect 19946 14592 21546 14648
rect 21602 14592 21607 14648
rect 19885 14590 21607 14592
rect 19885 14587 19951 14590
rect 21541 14587 21607 14590
rect 21950 14588 21956 14652
rect 22020 14650 22026 14652
rect 22185 14650 22251 14653
rect 22020 14648 22251 14650
rect 22020 14592 22190 14648
rect 22246 14592 22251 14648
rect 22020 14590 22251 14592
rect 22020 14588 22026 14590
rect 22185 14587 22251 14590
rect 22093 14514 22159 14517
rect 23105 14514 23171 14517
rect 22093 14512 23171 14514
rect 22093 14456 22098 14512
rect 22154 14456 23110 14512
rect 23166 14456 23171 14512
rect 22093 14454 23171 14456
rect 22093 14451 22159 14454
rect 23105 14451 23171 14454
rect 22461 14378 22527 14381
rect 26785 14378 26851 14381
rect 22461 14376 26851 14378
rect 22461 14320 22466 14376
rect 22522 14320 26790 14376
rect 26846 14320 26851 14376
rect 22461 14318 26851 14320
rect 22461 14315 22527 14318
rect 26785 14315 26851 14318
rect 22001 14242 22067 14245
rect 23473 14242 23539 14245
rect 22001 14240 23539 14242
rect 22001 14184 22006 14240
rect 22062 14184 23478 14240
rect 23534 14184 23539 14240
rect 22001 14182 23539 14184
rect 22001 14179 22067 14182
rect 23473 14179 23539 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 19333 13970 19399 13973
rect 20529 13970 20595 13973
rect 19333 13968 20595 13970
rect 19333 13912 19338 13968
rect 19394 13912 20534 13968
rect 20590 13912 20595 13968
rect 19333 13910 20595 13912
rect 19333 13907 19399 13910
rect 20529 13907 20595 13910
rect 18689 13834 18755 13837
rect 20345 13834 20411 13837
rect 18689 13832 20411 13834
rect 18689 13776 18694 13832
rect 18750 13776 20350 13832
rect 20406 13776 20411 13832
rect 18689 13774 20411 13776
rect 18689 13771 18755 13774
rect 20345 13771 20411 13774
rect 20989 13836 21055 13837
rect 20989 13832 21036 13836
rect 21100 13834 21106 13836
rect 20989 13776 20994 13832
rect 20989 13772 21036 13776
rect 21100 13774 21146 13834
rect 21100 13772 21106 13774
rect 20989 13771 21055 13772
rect 19149 13700 19215 13701
rect 19149 13696 19196 13700
rect 19260 13698 19266 13700
rect 24025 13698 24091 13701
rect 25681 13698 25747 13701
rect 19149 13640 19154 13696
rect 19149 13636 19196 13640
rect 19260 13638 19306 13698
rect 24025 13696 25747 13698
rect 24025 13640 24030 13696
rect 24086 13640 25686 13696
rect 25742 13640 25747 13696
rect 24025 13638 25747 13640
rect 19260 13636 19266 13638
rect 19149 13635 19215 13636
rect 24025 13635 24091 13638
rect 25681 13635 25747 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 20294 13500 20300 13564
rect 20364 13562 20370 13564
rect 20989 13562 21055 13565
rect 20364 13560 21055 13562
rect 20364 13504 20994 13560
rect 21050 13504 21055 13560
rect 20364 13502 21055 13504
rect 20364 13500 20370 13502
rect 20989 13499 21055 13502
rect 19517 13426 19583 13429
rect 20345 13426 20411 13429
rect 19517 13424 20411 13426
rect 19517 13368 19522 13424
rect 19578 13368 20350 13424
rect 20406 13368 20411 13424
rect 19517 13366 20411 13368
rect 19517 13363 19583 13366
rect 20345 13363 20411 13366
rect 13997 13290 14063 13293
rect 21725 13290 21791 13293
rect 13997 13288 21791 13290
rect 13997 13232 14002 13288
rect 14058 13232 21730 13288
rect 21786 13232 21791 13288
rect 13997 13230 21791 13232
rect 13997 13227 14063 13230
rect 21725 13227 21791 13230
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 14774 12820 14780 12884
rect 14844 12882 14850 12884
rect 15377 12882 15443 12885
rect 14844 12880 15443 12882
rect 14844 12824 15382 12880
rect 15438 12824 15443 12880
rect 14844 12822 15443 12824
rect 14844 12820 14850 12822
rect 15377 12819 15443 12822
rect 22185 12746 22251 12749
rect 24117 12746 24183 12749
rect 22185 12744 24183 12746
rect 22185 12688 22190 12744
rect 22246 12688 24122 12744
rect 24178 12688 24183 12744
rect 22185 12686 24183 12688
rect 22185 12683 22251 12686
rect 24117 12683 24183 12686
rect 22461 12610 22527 12613
rect 22737 12610 22803 12613
rect 22461 12608 22803 12610
rect 22461 12552 22466 12608
rect 22522 12552 22742 12608
rect 22798 12552 22803 12608
rect 22461 12550 22803 12552
rect 22461 12547 22527 12550
rect 22737 12547 22803 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 27981 12338 28047 12341
rect 28165 12338 28231 12341
rect 27981 12336 28231 12338
rect 27981 12280 27986 12336
rect 28042 12280 28170 12336
rect 28226 12280 28231 12336
rect 27981 12278 28231 12280
rect 27981 12275 28047 12278
rect 28165 12275 28231 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 20621 11794 20687 11797
rect 22829 11794 22895 11797
rect 20621 11792 22895 11794
rect 20621 11736 20626 11792
rect 20682 11736 22834 11792
rect 22890 11736 22895 11792
rect 20621 11734 22895 11736
rect 20621 11731 20687 11734
rect 22829 11731 22895 11734
rect 23105 11658 23171 11661
rect 26509 11658 26575 11661
rect 23105 11656 26575 11658
rect 23105 11600 23110 11656
rect 23166 11600 26514 11656
rect 26570 11600 26575 11656
rect 23105 11598 26575 11600
rect 23105 11595 23171 11598
rect 26509 11595 26575 11598
rect 20478 11460 20484 11524
rect 20548 11522 20554 11524
rect 20621 11522 20687 11525
rect 20548 11520 20687 11522
rect 20548 11464 20626 11520
rect 20682 11464 20687 11520
rect 20548 11462 20687 11464
rect 20548 11460 20554 11462
rect 20621 11459 20687 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 26325 11386 26391 11389
rect 19290 11384 26391 11386
rect 19290 11328 26330 11384
rect 26386 11328 26391 11384
rect 19290 11326 26391 11328
rect 16665 11250 16731 11253
rect 18505 11250 18571 11253
rect 16665 11248 18571 11250
rect 16665 11192 16670 11248
rect 16726 11192 18510 11248
rect 18566 11192 18571 11248
rect 16665 11190 18571 11192
rect 16665 11187 16731 11190
rect 18505 11187 18571 11190
rect 15101 11114 15167 11117
rect 19290 11114 19350 11326
rect 26325 11323 26391 11326
rect 23197 11250 23263 11253
rect 25957 11250 26023 11253
rect 23197 11248 26023 11250
rect 23197 11192 23202 11248
rect 23258 11192 25962 11248
rect 26018 11192 26023 11248
rect 23197 11190 26023 11192
rect 23197 11187 23263 11190
rect 25957 11187 26023 11190
rect 26734 11188 26740 11252
rect 26804 11250 26810 11252
rect 31477 11250 31543 11253
rect 26804 11248 31543 11250
rect 26804 11192 31482 11248
rect 31538 11192 31543 11248
rect 26804 11190 31543 11192
rect 26804 11188 26810 11190
rect 31477 11187 31543 11190
rect 15101 11112 19350 11114
rect 15101 11056 15106 11112
rect 15162 11056 19350 11112
rect 15101 11054 19350 11056
rect 25497 11114 25563 11117
rect 27521 11114 27587 11117
rect 25497 11112 27587 11114
rect 25497 11056 25502 11112
rect 25558 11056 27526 11112
rect 27582 11056 27587 11112
rect 25497 11054 27587 11056
rect 15101 11051 15167 11054
rect 25497 11051 25563 11054
rect 27521 11051 27587 11054
rect 16941 10978 17007 10981
rect 17861 10978 17927 10981
rect 16941 10976 17927 10978
rect 16941 10920 16946 10976
rect 17002 10920 17866 10976
rect 17922 10920 17927 10976
rect 16941 10918 17927 10920
rect 16941 10915 17007 10918
rect 17861 10915 17927 10918
rect 21081 10978 21147 10981
rect 21725 10978 21791 10981
rect 23565 10978 23631 10981
rect 21081 10976 23631 10978
rect 21081 10920 21086 10976
rect 21142 10920 21730 10976
rect 21786 10920 23570 10976
rect 23626 10920 23631 10976
rect 21081 10918 23631 10920
rect 21081 10915 21147 10918
rect 21725 10915 21791 10918
rect 23565 10915 23631 10918
rect 26049 10978 26115 10981
rect 26693 10978 26759 10981
rect 27797 10978 27863 10981
rect 26049 10976 27863 10978
rect 26049 10920 26054 10976
rect 26110 10920 26698 10976
rect 26754 10920 27802 10976
rect 27858 10920 27863 10976
rect 26049 10918 27863 10920
rect 26049 10915 26115 10918
rect 26693 10915 26759 10918
rect 27797 10915 27863 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 20662 10780 20668 10844
rect 20732 10842 20738 10844
rect 26877 10842 26943 10845
rect 20732 10840 26943 10842
rect 20732 10784 26882 10840
rect 26938 10784 26943 10840
rect 20732 10782 26943 10784
rect 20732 10780 20738 10782
rect 26877 10779 26943 10782
rect 19241 10708 19307 10709
rect 19190 10706 19196 10708
rect 19150 10646 19196 10706
rect 19260 10704 19307 10708
rect 19302 10648 19307 10704
rect 19190 10644 19196 10646
rect 19260 10644 19307 10648
rect 19241 10643 19307 10644
rect 23933 10706 23999 10709
rect 28717 10706 28783 10709
rect 23933 10704 28783 10706
rect 23933 10648 23938 10704
rect 23994 10648 28722 10704
rect 28778 10648 28783 10704
rect 23933 10646 28783 10648
rect 23933 10643 23999 10646
rect 28717 10643 28783 10646
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 22921 10298 22987 10301
rect 23381 10298 23447 10301
rect 22921 10296 23447 10298
rect 22921 10240 22926 10296
rect 22982 10240 23386 10296
rect 23442 10240 23447 10296
rect 22921 10238 23447 10240
rect 22921 10235 22987 10238
rect 23381 10235 23447 10238
rect 20253 10162 20319 10165
rect 22921 10162 22987 10165
rect 20253 10160 22987 10162
rect 20253 10104 20258 10160
rect 20314 10104 22926 10160
rect 22982 10104 22987 10160
rect 20253 10102 22987 10104
rect 20253 10099 20319 10102
rect 22921 10099 22987 10102
rect 20110 9964 20116 10028
rect 20180 10026 20186 10028
rect 21449 10026 21515 10029
rect 20180 10024 21515 10026
rect 20180 9968 21454 10024
rect 21510 9968 21515 10024
rect 20180 9966 21515 9968
rect 20180 9964 20186 9966
rect 21449 9963 21515 9966
rect 29545 9890 29611 9893
rect 30741 9890 30807 9893
rect 29545 9888 30807 9890
rect 29545 9832 29550 9888
rect 29606 9832 30746 9888
rect 30802 9832 30807 9888
rect 29545 9830 30807 9832
rect 29545 9827 29611 9830
rect 30741 9827 30807 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 10777 9618 10843 9621
rect 13261 9618 13327 9621
rect 17493 9620 17559 9621
rect 17493 9618 17540 9620
rect 10777 9616 13327 9618
rect 10777 9560 10782 9616
rect 10838 9560 13266 9616
rect 13322 9560 13327 9616
rect 10777 9558 13327 9560
rect 17448 9616 17540 9618
rect 17448 9560 17498 9616
rect 17448 9558 17540 9560
rect 10777 9555 10843 9558
rect 13261 9555 13327 9558
rect 17493 9556 17540 9558
rect 17604 9556 17610 9620
rect 21817 9618 21883 9621
rect 22369 9618 22435 9621
rect 21817 9616 22435 9618
rect 21817 9560 21822 9616
rect 21878 9560 22374 9616
rect 22430 9560 22435 9616
rect 21817 9558 22435 9560
rect 17493 9555 17559 9556
rect 21817 9555 21883 9558
rect 22369 9555 22435 9558
rect 22645 9618 22711 9621
rect 24025 9618 24091 9621
rect 22645 9616 24091 9618
rect 22645 9560 22650 9616
rect 22706 9560 24030 9616
rect 24086 9560 24091 9616
rect 22645 9558 24091 9560
rect 22645 9555 22711 9558
rect 24025 9555 24091 9558
rect 24669 9618 24735 9621
rect 25681 9618 25747 9621
rect 24669 9616 25747 9618
rect 24669 9560 24674 9616
rect 24730 9560 25686 9616
rect 25742 9560 25747 9616
rect 24669 9558 25747 9560
rect 24669 9555 24735 9558
rect 25681 9555 25747 9558
rect 16941 9482 17007 9485
rect 19057 9482 19123 9485
rect 16941 9480 19123 9482
rect 16941 9424 16946 9480
rect 17002 9424 19062 9480
rect 19118 9424 19123 9480
rect 16941 9422 19123 9424
rect 16941 9419 17007 9422
rect 19057 9419 19123 9422
rect 20110 9420 20116 9484
rect 20180 9482 20186 9484
rect 26509 9482 26575 9485
rect 20180 9480 26575 9482
rect 20180 9424 26514 9480
rect 26570 9424 26575 9480
rect 20180 9422 26575 9424
rect 20180 9420 20186 9422
rect 26509 9419 26575 9422
rect 27705 9482 27771 9485
rect 30557 9482 30623 9485
rect 27705 9480 30623 9482
rect 27705 9424 27710 9480
rect 27766 9424 30562 9480
rect 30618 9424 30623 9480
rect 27705 9422 30623 9424
rect 27705 9419 27771 9422
rect 30557 9419 30623 9422
rect 17217 9346 17283 9349
rect 19977 9346 20043 9349
rect 17217 9344 20043 9346
rect 17217 9288 17222 9344
rect 17278 9288 19982 9344
rect 20038 9288 20043 9344
rect 17217 9286 20043 9288
rect 17217 9283 17283 9286
rect 19977 9283 20043 9286
rect 22093 9346 22159 9349
rect 27889 9346 27955 9349
rect 22093 9344 27955 9346
rect 22093 9288 22098 9344
rect 22154 9288 27894 9344
rect 27950 9288 27955 9344
rect 22093 9286 27955 9288
rect 22093 9283 22159 9286
rect 27889 9283 27955 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 16849 9210 16915 9213
rect 18597 9210 18663 9213
rect 16849 9208 18663 9210
rect 16849 9152 16854 9208
rect 16910 9152 18602 9208
rect 18658 9152 18663 9208
rect 16849 9150 18663 9152
rect 16849 9147 16915 9150
rect 18597 9147 18663 9150
rect 19517 9210 19583 9213
rect 27613 9210 27679 9213
rect 19517 9208 27679 9210
rect 19517 9152 19522 9208
rect 19578 9152 27618 9208
rect 27674 9152 27679 9208
rect 19517 9150 27679 9152
rect 19517 9147 19583 9150
rect 27613 9147 27679 9150
rect 3969 9074 4035 9077
rect 7465 9074 7531 9077
rect 3969 9072 7531 9074
rect 3969 9016 3974 9072
rect 4030 9016 7470 9072
rect 7526 9016 7531 9072
rect 3969 9014 7531 9016
rect 3969 9011 4035 9014
rect 7465 9011 7531 9014
rect 13445 9074 13511 9077
rect 18873 9074 18939 9077
rect 13445 9072 18939 9074
rect 13445 9016 13450 9072
rect 13506 9016 18878 9072
rect 18934 9016 18939 9072
rect 13445 9014 18939 9016
rect 13445 9011 13511 9014
rect 18873 9011 18939 9014
rect 22001 9074 22067 9077
rect 22645 9074 22711 9077
rect 22001 9072 22711 9074
rect 22001 9016 22006 9072
rect 22062 9016 22650 9072
rect 22706 9016 22711 9072
rect 22001 9014 22711 9016
rect 22001 9011 22067 9014
rect 22645 9011 22711 9014
rect 27521 9074 27587 9077
rect 30649 9074 30715 9077
rect 27521 9072 30715 9074
rect 27521 9016 27526 9072
rect 27582 9016 30654 9072
rect 30710 9016 30715 9072
rect 27521 9014 30715 9016
rect 27521 9011 27587 9014
rect 30649 9011 30715 9014
rect 10041 8938 10107 8941
rect 15377 8938 15443 8941
rect 10041 8936 15443 8938
rect 10041 8880 10046 8936
rect 10102 8880 15382 8936
rect 15438 8880 15443 8936
rect 10041 8878 15443 8880
rect 10041 8875 10107 8878
rect 15377 8875 15443 8878
rect 21817 8936 21883 8941
rect 21817 8880 21822 8936
rect 21878 8880 21883 8936
rect 21817 8875 21883 8880
rect 27061 8938 27127 8941
rect 28533 8938 28599 8941
rect 27061 8936 28599 8938
rect 27061 8880 27066 8936
rect 27122 8880 28538 8936
rect 28594 8880 28599 8936
rect 27061 8878 28599 8880
rect 27061 8875 27127 8878
rect 28533 8875 28599 8878
rect 4153 8802 4219 8805
rect 10409 8802 10475 8805
rect 4153 8800 10475 8802
rect 4153 8744 4158 8800
rect 4214 8744 10414 8800
rect 10470 8744 10475 8800
rect 4153 8742 10475 8744
rect 4153 8739 4219 8742
rect 10409 8739 10475 8742
rect 12525 8802 12591 8805
rect 17534 8802 17540 8804
rect 12525 8800 17540 8802
rect 12525 8744 12530 8800
rect 12586 8744 17540 8800
rect 12525 8742 17540 8744
rect 12525 8739 12591 8742
rect 17534 8740 17540 8742
rect 17604 8802 17610 8804
rect 18321 8802 18387 8805
rect 17604 8800 18387 8802
rect 17604 8744 18326 8800
rect 18382 8744 18387 8800
rect 17604 8742 18387 8744
rect 17604 8740 17610 8742
rect 18321 8739 18387 8742
rect 20846 8740 20852 8804
rect 20916 8802 20922 8804
rect 20989 8802 21055 8805
rect 20916 8800 21055 8802
rect 20916 8744 20994 8800
rect 21050 8744 21055 8800
rect 20916 8742 21055 8744
rect 21820 8802 21880 8875
rect 29085 8802 29151 8805
rect 21820 8800 29151 8802
rect 21820 8744 29090 8800
rect 29146 8744 29151 8800
rect 21820 8742 29151 8744
rect 20916 8740 20922 8742
rect 20989 8739 21055 8742
rect 29085 8739 29151 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 4061 8666 4127 8669
rect 9305 8666 9371 8669
rect 4061 8664 9371 8666
rect 4061 8608 4066 8664
rect 4122 8608 9310 8664
rect 9366 8608 9371 8664
rect 4061 8606 9371 8608
rect 4061 8603 4127 8606
rect 9305 8603 9371 8606
rect 18413 8666 18479 8669
rect 19425 8666 19491 8669
rect 18413 8664 19491 8666
rect 18413 8608 18418 8664
rect 18474 8608 19430 8664
rect 19486 8608 19491 8664
rect 18413 8606 19491 8608
rect 18413 8603 18479 8606
rect 19425 8603 19491 8606
rect 20253 8666 20319 8669
rect 20805 8666 20871 8669
rect 20253 8664 20871 8666
rect 20253 8608 20258 8664
rect 20314 8608 20810 8664
rect 20866 8608 20871 8664
rect 20253 8606 20871 8608
rect 20253 8603 20319 8606
rect 20805 8603 20871 8606
rect 25037 8666 25103 8669
rect 28165 8666 28231 8669
rect 25037 8664 28231 8666
rect 25037 8608 25042 8664
rect 25098 8608 28170 8664
rect 28226 8608 28231 8664
rect 25037 8606 28231 8608
rect 25037 8603 25103 8606
rect 28165 8603 28231 8606
rect 3233 8530 3299 8533
rect 6913 8530 6979 8533
rect 3233 8528 6979 8530
rect 3233 8472 3238 8528
rect 3294 8472 6918 8528
rect 6974 8472 6979 8528
rect 3233 8470 6979 8472
rect 3233 8467 3299 8470
rect 6913 8467 6979 8470
rect 19190 8468 19196 8532
rect 19260 8530 19266 8532
rect 19977 8530 20043 8533
rect 19260 8528 20043 8530
rect 19260 8472 19982 8528
rect 20038 8472 20043 8528
rect 19260 8470 20043 8472
rect 19260 8468 19266 8470
rect 19977 8467 20043 8470
rect 3601 8394 3667 8397
rect 7005 8394 7071 8397
rect 3601 8392 7071 8394
rect 3601 8336 3606 8392
rect 3662 8336 7010 8392
rect 7066 8336 7071 8392
rect 3601 8334 7071 8336
rect 3601 8331 3667 8334
rect 7005 8331 7071 8334
rect 20437 8394 20503 8397
rect 22001 8394 22067 8397
rect 20437 8392 22067 8394
rect 20437 8336 20442 8392
rect 20498 8336 22006 8392
rect 22062 8336 22067 8392
rect 20437 8334 22067 8336
rect 20437 8331 20503 8334
rect 22001 8331 22067 8334
rect 23013 8394 23079 8397
rect 23289 8394 23355 8397
rect 23013 8392 23355 8394
rect 23013 8336 23018 8392
rect 23074 8336 23294 8392
rect 23350 8336 23355 8392
rect 23013 8334 23355 8336
rect 23013 8331 23079 8334
rect 23289 8331 23355 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 5073 8122 5139 8125
rect 5993 8122 6059 8125
rect 5073 8120 6059 8122
rect 5073 8064 5078 8120
rect 5134 8064 5998 8120
rect 6054 8064 6059 8120
rect 5073 8062 6059 8064
rect 5073 8059 5139 8062
rect 5993 8059 6059 8062
rect 4521 7850 4587 7853
rect 9673 7850 9739 7853
rect 4521 7848 9739 7850
rect 4521 7792 4526 7848
rect 4582 7792 9678 7848
rect 9734 7792 9739 7848
rect 4521 7790 9739 7792
rect 4521 7787 4587 7790
rect 9673 7787 9739 7790
rect 2313 7714 2379 7717
rect 5349 7714 5415 7717
rect 2313 7712 5415 7714
rect 2313 7656 2318 7712
rect 2374 7656 5354 7712
rect 5410 7656 5415 7712
rect 2313 7654 5415 7656
rect 2313 7651 2379 7654
rect 5349 7651 5415 7654
rect 22921 7714 22987 7717
rect 27429 7714 27495 7717
rect 22921 7712 27495 7714
rect 22921 7656 22926 7712
rect 22982 7656 27434 7712
rect 27490 7656 27495 7712
rect 22921 7654 27495 7656
rect 22921 7651 22987 7654
rect 27429 7651 27495 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3693 7578 3759 7581
rect 7833 7578 7899 7581
rect 3693 7576 7899 7578
rect 3693 7520 3698 7576
rect 3754 7520 7838 7576
rect 7894 7520 7899 7576
rect 3693 7518 7899 7520
rect 3693 7515 3759 7518
rect 7833 7515 7899 7518
rect 25814 7516 25820 7580
rect 25884 7578 25890 7580
rect 31937 7578 32003 7581
rect 25884 7576 32003 7578
rect 25884 7520 31942 7576
rect 31998 7520 32003 7576
rect 25884 7518 32003 7520
rect 25884 7516 25890 7518
rect 31937 7515 32003 7518
rect 3233 7442 3299 7445
rect 11513 7442 11579 7445
rect 3233 7440 11579 7442
rect 3233 7384 3238 7440
rect 3294 7384 11518 7440
rect 11574 7384 11579 7440
rect 3233 7382 11579 7384
rect 3233 7379 3299 7382
rect 11513 7379 11579 7382
rect 20437 7442 20503 7445
rect 28257 7442 28323 7445
rect 20437 7440 28323 7442
rect 20437 7384 20442 7440
rect 20498 7384 28262 7440
rect 28318 7384 28323 7440
rect 20437 7382 28323 7384
rect 20437 7379 20503 7382
rect 28257 7379 28323 7382
rect 4429 7306 4495 7309
rect 9765 7306 9831 7309
rect 4429 7304 9831 7306
rect 4429 7248 4434 7304
rect 4490 7248 9770 7304
rect 9826 7248 9831 7304
rect 4429 7246 9831 7248
rect 4429 7243 4495 7246
rect 9765 7243 9831 7246
rect 13629 7306 13695 7309
rect 15009 7306 15075 7309
rect 15561 7306 15627 7309
rect 13629 7304 15627 7306
rect 13629 7248 13634 7304
rect 13690 7248 15014 7304
rect 15070 7248 15566 7304
rect 15622 7248 15627 7304
rect 13629 7246 15627 7248
rect 13629 7243 13695 7246
rect 15009 7243 15075 7246
rect 15561 7243 15627 7246
rect 23289 7306 23355 7309
rect 27981 7306 28047 7309
rect 23289 7304 28047 7306
rect 23289 7248 23294 7304
rect 23350 7248 27986 7304
rect 28042 7248 28047 7304
rect 23289 7246 28047 7248
rect 23289 7243 23355 7246
rect 27981 7243 28047 7246
rect 4889 7170 4955 7173
rect 8293 7170 8359 7173
rect 4889 7168 8359 7170
rect 4889 7112 4894 7168
rect 4950 7112 8298 7168
rect 8354 7112 8359 7168
rect 4889 7110 8359 7112
rect 4889 7107 4955 7110
rect 8293 7107 8359 7110
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 5349 6898 5415 6901
rect 9489 6898 9555 6901
rect 5349 6896 9555 6898
rect 5349 6840 5354 6896
rect 5410 6840 9494 6896
rect 9550 6840 9555 6896
rect 5349 6838 9555 6840
rect 5349 6835 5415 6838
rect 9489 6835 9555 6838
rect 15377 6898 15443 6901
rect 21030 6898 21036 6900
rect 15377 6896 21036 6898
rect 15377 6840 15382 6896
rect 15438 6840 21036 6896
rect 15377 6838 21036 6840
rect 15377 6835 15443 6838
rect 21030 6836 21036 6838
rect 21100 6836 21106 6900
rect 28022 6836 28028 6900
rect 28092 6898 28098 6900
rect 31293 6898 31359 6901
rect 28092 6896 31359 6898
rect 28092 6840 31298 6896
rect 31354 6840 31359 6896
rect 28092 6838 31359 6840
rect 28092 6836 28098 6838
rect 31293 6835 31359 6838
rect 31477 6898 31543 6901
rect 31753 6898 31819 6901
rect 31477 6896 31819 6898
rect 31477 6840 31482 6896
rect 31538 6840 31758 6896
rect 31814 6840 31819 6896
rect 31477 6838 31819 6840
rect 31477 6835 31543 6838
rect 31753 6835 31819 6838
rect 17585 6762 17651 6765
rect 23238 6762 23244 6764
rect 17585 6760 23244 6762
rect 17585 6704 17590 6760
rect 17646 6704 23244 6760
rect 17585 6702 23244 6704
rect 17585 6699 17651 6702
rect 23238 6700 23244 6702
rect 23308 6700 23314 6764
rect 29913 6762 29979 6765
rect 28950 6760 29979 6762
rect 28950 6704 29918 6760
rect 29974 6704 29979 6760
rect 28950 6702 29979 6704
rect 20989 6626 21055 6629
rect 28950 6626 29010 6702
rect 29913 6699 29979 6702
rect 20989 6624 29010 6626
rect 20989 6568 20994 6624
rect 21050 6568 29010 6624
rect 20989 6566 29010 6568
rect 20989 6563 21055 6566
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 1669 6490 1735 6493
rect 6637 6490 6703 6493
rect 1669 6488 6703 6490
rect 1669 6432 1674 6488
rect 1730 6432 6642 6488
rect 6698 6432 6703 6488
rect 1669 6430 6703 6432
rect 1669 6427 1735 6430
rect 6637 6427 6703 6430
rect 6913 6490 6979 6493
rect 8937 6490 9003 6493
rect 6913 6488 9003 6490
rect 6913 6432 6918 6488
rect 6974 6432 8942 6488
rect 8998 6432 9003 6488
rect 6913 6430 9003 6432
rect 6913 6427 6979 6430
rect 8937 6427 9003 6430
rect 3693 6354 3759 6357
rect 9673 6354 9739 6357
rect 3693 6352 9739 6354
rect 3693 6296 3698 6352
rect 3754 6296 9678 6352
rect 9734 6296 9739 6352
rect 3693 6294 9739 6296
rect 3693 6291 3759 6294
rect 9673 6291 9739 6294
rect 11881 6354 11947 6357
rect 12617 6354 12683 6357
rect 11881 6352 12683 6354
rect 11881 6296 11886 6352
rect 11942 6296 12622 6352
rect 12678 6296 12683 6352
rect 11881 6294 12683 6296
rect 11881 6291 11947 6294
rect 12617 6291 12683 6294
rect 19885 6354 19951 6357
rect 20989 6354 21055 6357
rect 19885 6352 21055 6354
rect 19885 6296 19890 6352
rect 19946 6296 20994 6352
rect 21050 6296 21055 6352
rect 19885 6294 21055 6296
rect 19885 6291 19951 6294
rect 20989 6291 21055 6294
rect 22369 6354 22435 6357
rect 24301 6354 24367 6357
rect 22369 6352 24367 6354
rect 22369 6296 22374 6352
rect 22430 6296 24306 6352
rect 24362 6296 24367 6352
rect 22369 6294 24367 6296
rect 22369 6291 22435 6294
rect 24301 6291 24367 6294
rect 3693 6218 3759 6221
rect 8385 6218 8451 6221
rect 3693 6216 8451 6218
rect 3693 6160 3698 6216
rect 3754 6160 8390 6216
rect 8446 6160 8451 6216
rect 3693 6158 8451 6160
rect 3693 6155 3759 6158
rect 8385 6155 8451 6158
rect 10317 6218 10383 6221
rect 16297 6218 16363 6221
rect 10317 6216 16363 6218
rect 10317 6160 10322 6216
rect 10378 6160 16302 6216
rect 16358 6160 16363 6216
rect 10317 6158 16363 6160
rect 10317 6155 10383 6158
rect 16297 6155 16363 6158
rect 20529 6218 20595 6221
rect 26734 6218 26740 6220
rect 20529 6216 26740 6218
rect 20529 6160 20534 6216
rect 20590 6160 26740 6216
rect 20529 6158 26740 6160
rect 20529 6155 20595 6158
rect 26734 6156 26740 6158
rect 26804 6156 26810 6220
rect 5073 6082 5139 6085
rect 8293 6082 8359 6085
rect 5073 6080 8359 6082
rect 5073 6024 5078 6080
rect 5134 6024 8298 6080
rect 8354 6024 8359 6080
rect 5073 6022 8359 6024
rect 5073 6019 5139 6022
rect 8293 6019 8359 6022
rect 23473 6082 23539 6085
rect 25129 6082 25195 6085
rect 23473 6080 25195 6082
rect 23473 6024 23478 6080
rect 23534 6024 25134 6080
rect 25190 6024 25195 6080
rect 23473 6022 25195 6024
rect 23473 6019 23539 6022
rect 25129 6019 25195 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 23381 5946 23447 5949
rect 27981 5946 28047 5949
rect 23381 5944 28047 5946
rect 23381 5888 23386 5944
rect 23442 5888 27986 5944
rect 28042 5888 28047 5944
rect 23381 5886 28047 5888
rect 23381 5883 23447 5886
rect 27981 5883 28047 5886
rect 4981 5810 5047 5813
rect 8661 5810 8727 5813
rect 4981 5808 8727 5810
rect 4981 5752 4986 5808
rect 5042 5752 8666 5808
rect 8722 5752 8727 5808
rect 4981 5750 8727 5752
rect 4981 5747 5047 5750
rect 8661 5747 8727 5750
rect 25773 5810 25839 5813
rect 27429 5810 27495 5813
rect 25773 5808 27495 5810
rect 25773 5752 25778 5808
rect 25834 5752 27434 5808
rect 27490 5752 27495 5808
rect 25773 5750 27495 5752
rect 25773 5747 25839 5750
rect 27429 5747 27495 5750
rect 3693 5674 3759 5677
rect 10869 5674 10935 5677
rect 3693 5672 10935 5674
rect 3693 5616 3698 5672
rect 3754 5616 10874 5672
rect 10930 5616 10935 5672
rect 3693 5614 10935 5616
rect 3693 5611 3759 5614
rect 10869 5611 10935 5614
rect 26877 5674 26943 5677
rect 28073 5674 28139 5677
rect 26877 5672 28139 5674
rect 26877 5616 26882 5672
rect 26938 5616 28078 5672
rect 28134 5616 28139 5672
rect 26877 5614 28139 5616
rect 26877 5611 26943 5614
rect 28073 5611 28139 5614
rect 2497 5538 2563 5541
rect 7005 5538 7071 5541
rect 2497 5536 7071 5538
rect 2497 5480 2502 5536
rect 2558 5480 7010 5536
rect 7066 5480 7071 5536
rect 2497 5478 7071 5480
rect 2497 5475 2563 5478
rect 7005 5475 7071 5478
rect 7465 5538 7531 5541
rect 10225 5538 10291 5541
rect 7465 5536 10291 5538
rect 7465 5480 7470 5536
rect 7526 5480 10230 5536
rect 10286 5480 10291 5536
rect 7465 5478 10291 5480
rect 7465 5475 7531 5478
rect 10225 5475 10291 5478
rect 10961 5538 11027 5541
rect 12617 5538 12683 5541
rect 10961 5536 12683 5538
rect 10961 5480 10966 5536
rect 11022 5480 12622 5536
rect 12678 5480 12683 5536
rect 10961 5478 12683 5480
rect 10961 5475 11027 5478
rect 12617 5475 12683 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 3141 5402 3207 5405
rect 11329 5402 11395 5405
rect 3141 5400 11395 5402
rect 3141 5344 3146 5400
rect 3202 5344 11334 5400
rect 11390 5344 11395 5400
rect 3141 5342 11395 5344
rect 3141 5339 3207 5342
rect 11329 5339 11395 5342
rect 3417 5266 3483 5269
rect 4889 5266 4955 5269
rect 3417 5264 4955 5266
rect 3417 5208 3422 5264
rect 3478 5208 4894 5264
rect 4950 5208 4955 5264
rect 3417 5206 4955 5208
rect 3417 5203 3483 5206
rect 4889 5203 4955 5206
rect 1853 5130 1919 5133
rect 11421 5130 11487 5133
rect 1853 5128 11487 5130
rect 1853 5072 1858 5128
rect 1914 5072 11426 5128
rect 11482 5072 11487 5128
rect 1853 5070 11487 5072
rect 1853 5067 1919 5070
rect 11421 5067 11487 5070
rect 9765 4994 9831 4997
rect 15469 4994 15535 4997
rect 9765 4992 15535 4994
rect 9765 4936 9770 4992
rect 9826 4936 15474 4992
rect 15530 4936 15535 4992
rect 9765 4934 15535 4936
rect 9765 4931 9831 4934
rect 15469 4931 15535 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 10409 4858 10475 4861
rect 10961 4858 11027 4861
rect 10409 4856 11027 4858
rect 10409 4800 10414 4856
rect 10470 4800 10966 4856
rect 11022 4800 11027 4856
rect 10409 4798 11027 4800
rect 10409 4795 10475 4798
rect 10961 4795 11027 4798
rect 3233 4722 3299 4725
rect 9857 4722 9923 4725
rect 3233 4720 9923 4722
rect 3233 4664 3238 4720
rect 3294 4664 9862 4720
rect 9918 4664 9923 4720
rect 3233 4662 9923 4664
rect 3233 4659 3299 4662
rect 9857 4659 9923 4662
rect 3785 4586 3851 4589
rect 6361 4586 6427 4589
rect 3785 4584 6427 4586
rect 3785 4528 3790 4584
rect 3846 4528 6366 4584
rect 6422 4528 6427 4584
rect 3785 4526 6427 4528
rect 3785 4523 3851 4526
rect 6361 4523 6427 4526
rect 3325 4450 3391 4453
rect 11973 4450 12039 4453
rect 3325 4448 12039 4450
rect 3325 4392 3330 4448
rect 3386 4392 11978 4448
rect 12034 4392 12039 4448
rect 3325 4390 12039 4392
rect 3325 4387 3391 4390
rect 11973 4387 12039 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 11053 4314 11119 4317
rect 3006 4312 11119 4314
rect 3006 4256 11058 4312
rect 11114 4256 11119 4312
rect 3006 4254 11119 4256
rect 2865 4178 2931 4181
rect 3006 4178 3066 4254
rect 11053 4251 11119 4254
rect 11513 4314 11579 4317
rect 11973 4314 12039 4317
rect 11513 4312 12039 4314
rect 11513 4256 11518 4312
rect 11574 4256 11978 4312
rect 12034 4256 12039 4312
rect 11513 4254 12039 4256
rect 11513 4251 11579 4254
rect 11973 4251 12039 4254
rect 2865 4176 3066 4178
rect 2865 4120 2870 4176
rect 2926 4120 3066 4176
rect 2865 4118 3066 4120
rect 3325 4178 3391 4181
rect 8937 4178 9003 4181
rect 3325 4176 9003 4178
rect 3325 4120 3330 4176
rect 3386 4120 8942 4176
rect 8998 4120 9003 4176
rect 3325 4118 9003 4120
rect 2865 4115 2931 4118
rect 3325 4115 3391 4118
rect 8937 4115 9003 4118
rect 9673 4176 9739 4181
rect 9673 4120 9678 4176
rect 9734 4120 9739 4176
rect 9673 4115 9739 4120
rect 14181 4178 14247 4181
rect 16665 4178 16731 4181
rect 14181 4176 16731 4178
rect 14181 4120 14186 4176
rect 14242 4120 16670 4176
rect 16726 4120 16731 4176
rect 14181 4118 16731 4120
rect 14181 4115 14247 4118
rect 16665 4115 16731 4118
rect 19609 4178 19675 4181
rect 20713 4178 20779 4181
rect 19609 4176 20779 4178
rect 19609 4120 19614 4176
rect 19670 4120 20718 4176
rect 20774 4120 20779 4176
rect 19609 4118 20779 4120
rect 19609 4115 19675 4118
rect 20713 4115 20779 4118
rect 28165 4178 28231 4181
rect 28809 4178 28875 4181
rect 28165 4176 28875 4178
rect 28165 4120 28170 4176
rect 28226 4120 28814 4176
rect 28870 4120 28875 4176
rect 28165 4118 28875 4120
rect 28165 4115 28231 4118
rect 28809 4115 28875 4118
rect 3601 4042 3667 4045
rect 9676 4042 9736 4115
rect 12709 4042 12775 4045
rect 3601 4040 7666 4042
rect 3601 3984 3606 4040
rect 3662 3984 7666 4040
rect 3601 3982 7666 3984
rect 9676 4040 12775 4042
rect 9676 3984 12714 4040
rect 12770 3984 12775 4040
rect 9676 3982 12775 3984
rect 3601 3979 3667 3982
rect 4889 3906 4955 3909
rect 5901 3906 5967 3909
rect 4889 3904 5967 3906
rect 4889 3848 4894 3904
rect 4950 3848 5906 3904
rect 5962 3848 5967 3904
rect 4889 3846 5967 3848
rect 7606 3906 7666 3982
rect 12709 3979 12775 3982
rect 14641 4042 14707 4045
rect 14774 4042 14780 4044
rect 14641 4040 14780 4042
rect 14641 3984 14646 4040
rect 14702 3984 14780 4040
rect 14641 3982 14780 3984
rect 14641 3979 14707 3982
rect 14774 3980 14780 3982
rect 14844 3980 14850 4044
rect 19149 4042 19215 4045
rect 20345 4044 20411 4045
rect 20110 4042 20116 4044
rect 19149 4040 20116 4042
rect 19149 3984 19154 4040
rect 19210 3984 20116 4040
rect 19149 3982 20116 3984
rect 19149 3979 19215 3982
rect 20110 3980 20116 3982
rect 20180 3980 20186 4044
rect 20294 3980 20300 4044
rect 20364 4042 20411 4044
rect 20989 4042 21055 4045
rect 28022 4042 28028 4044
rect 20364 4040 20456 4042
rect 20406 3984 20456 4040
rect 20364 3982 20456 3984
rect 20989 4040 28028 4042
rect 20989 3984 20994 4040
rect 21050 3984 28028 4040
rect 20989 3982 28028 3984
rect 20364 3980 20411 3982
rect 20345 3979 20411 3980
rect 20989 3979 21055 3982
rect 28022 3980 28028 3982
rect 28092 3980 28098 4044
rect 8293 3906 8359 3909
rect 7606 3904 8359 3906
rect 7606 3848 8298 3904
rect 8354 3848 8359 3904
rect 7606 3846 8359 3848
rect 4889 3843 4955 3846
rect 5901 3843 5967 3846
rect 8293 3843 8359 3846
rect 11973 3906 12039 3909
rect 17033 3906 17099 3909
rect 11973 3904 17099 3906
rect 11973 3848 11978 3904
rect 12034 3848 17038 3904
rect 17094 3848 17099 3904
rect 11973 3846 17099 3848
rect 11973 3843 12039 3846
rect 17033 3843 17099 3846
rect 19517 3906 19583 3909
rect 23289 3906 23355 3909
rect 19517 3904 23355 3906
rect 19517 3848 19522 3904
rect 19578 3848 23294 3904
rect 23350 3848 23355 3904
rect 19517 3846 23355 3848
rect 19517 3843 19583 3846
rect 23289 3843 23355 3846
rect 25681 3906 25747 3909
rect 25814 3906 25820 3908
rect 25681 3904 25820 3906
rect 25681 3848 25686 3904
rect 25742 3848 25820 3904
rect 25681 3846 25820 3848
rect 25681 3843 25747 3846
rect 25814 3844 25820 3846
rect 25884 3844 25890 3908
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 5533 3770 5599 3773
rect 6177 3770 6243 3773
rect 5533 3768 6243 3770
rect 5533 3712 5538 3768
rect 5594 3712 6182 3768
rect 6238 3712 6243 3768
rect 5533 3710 6243 3712
rect 5533 3707 5599 3710
rect 6177 3707 6243 3710
rect 12249 3770 12315 3773
rect 16757 3770 16823 3773
rect 12249 3768 16823 3770
rect 12249 3712 12254 3768
rect 12310 3712 16762 3768
rect 16818 3712 16823 3768
rect 12249 3710 16823 3712
rect 12249 3707 12315 3710
rect 16757 3707 16823 3710
rect 19793 3770 19859 3773
rect 23473 3770 23539 3773
rect 19793 3768 23539 3770
rect 19793 3712 19798 3768
rect 19854 3712 23478 3768
rect 23534 3712 23539 3768
rect 19793 3710 23539 3712
rect 19793 3707 19859 3710
rect 23473 3707 23539 3710
rect 3417 3634 3483 3637
rect 8385 3634 8451 3637
rect 3417 3632 8451 3634
rect 3417 3576 3422 3632
rect 3478 3576 8390 3632
rect 8446 3576 8451 3632
rect 3417 3574 8451 3576
rect 3417 3571 3483 3574
rect 8385 3571 8451 3574
rect 10593 3634 10659 3637
rect 12341 3634 12407 3637
rect 10593 3632 12407 3634
rect 10593 3576 10598 3632
rect 10654 3576 12346 3632
rect 12402 3576 12407 3632
rect 10593 3574 12407 3576
rect 10593 3571 10659 3574
rect 12341 3571 12407 3574
rect 14273 3634 14339 3637
rect 14825 3634 14891 3637
rect 14273 3632 14891 3634
rect 14273 3576 14278 3632
rect 14334 3576 14830 3632
rect 14886 3576 14891 3632
rect 14273 3574 14891 3576
rect 14273 3571 14339 3574
rect 14825 3571 14891 3574
rect 18229 3634 18295 3637
rect 19333 3634 19399 3637
rect 18229 3632 19399 3634
rect 18229 3576 18234 3632
rect 18290 3576 19338 3632
rect 19394 3576 19399 3632
rect 18229 3574 19399 3576
rect 18229 3571 18295 3574
rect 19333 3571 19399 3574
rect 20253 3634 20319 3637
rect 20805 3634 20871 3637
rect 20253 3632 20871 3634
rect 20253 3576 20258 3632
rect 20314 3576 20810 3632
rect 20866 3576 20871 3632
rect 20253 3574 20871 3576
rect 20253 3571 20319 3574
rect 20805 3571 20871 3574
rect 3785 3498 3851 3501
rect 13169 3498 13235 3501
rect 3785 3496 13235 3498
rect 3785 3440 3790 3496
rect 3846 3440 13174 3496
rect 13230 3440 13235 3496
rect 3785 3438 13235 3440
rect 3785 3435 3851 3438
rect 13169 3435 13235 3438
rect 19425 3498 19491 3501
rect 19425 3496 20040 3498
rect 19425 3440 19430 3496
rect 19486 3440 20040 3496
rect 19425 3438 20040 3440
rect 19425 3435 19491 3438
rect 197 3362 263 3365
rect 19374 3362 19380 3364
rect 197 3360 19380 3362
rect 197 3304 202 3360
rect 258 3304 19380 3360
rect 197 3302 19380 3304
rect 197 3299 263 3302
rect 19374 3300 19380 3302
rect 19444 3300 19450 3364
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 3141 3226 3207 3229
rect 8569 3226 8635 3229
rect 3141 3224 8635 3226
rect 3141 3168 3146 3224
rect 3202 3168 8574 3224
rect 8630 3168 8635 3224
rect 3141 3166 8635 3168
rect 3141 3163 3207 3166
rect 8569 3163 8635 3166
rect 1669 3090 1735 3093
rect 7189 3090 7255 3093
rect 1669 3088 7255 3090
rect 1669 3032 1674 3088
rect 1730 3032 7194 3088
rect 7250 3032 7255 3088
rect 1669 3030 7255 3032
rect 1669 3027 1735 3030
rect 7189 3027 7255 3030
rect 7465 3090 7531 3093
rect 9121 3090 9187 3093
rect 7465 3088 9187 3090
rect 7465 3032 7470 3088
rect 7526 3032 9126 3088
rect 9182 3032 9187 3088
rect 7465 3030 9187 3032
rect 7465 3027 7531 3030
rect 9121 3027 9187 3030
rect 3141 2954 3207 2957
rect 9305 2954 9371 2957
rect 3141 2952 9371 2954
rect 3141 2896 3146 2952
rect 3202 2896 9310 2952
rect 9366 2896 9371 2952
rect 3141 2894 9371 2896
rect 3141 2891 3207 2894
rect 9305 2891 9371 2894
rect 19425 2954 19491 2957
rect 19980 2954 20040 3438
rect 19425 2952 20040 2954
rect 19425 2896 19430 2952
rect 19486 2896 20040 2952
rect 19425 2894 20040 2896
rect 20529 2954 20595 2957
rect 20662 2954 20668 2956
rect 20529 2952 20668 2954
rect 20529 2896 20534 2952
rect 20590 2896 20668 2952
rect 20529 2894 20668 2896
rect 19425 2891 19491 2894
rect 20529 2891 20595 2894
rect 20662 2892 20668 2894
rect 20732 2892 20738 2956
rect 19793 2818 19859 2821
rect 28717 2818 28783 2821
rect 19793 2816 28783 2818
rect 19793 2760 19798 2816
rect 19854 2760 28722 2816
rect 28778 2760 28783 2816
rect 19793 2758 28783 2760
rect 19793 2755 19859 2758
rect 28717 2755 28783 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 19517 2546 19583 2549
rect 20294 2546 20300 2548
rect 19517 2544 20300 2546
rect 19517 2488 19522 2544
rect 19578 2488 20300 2544
rect 19517 2486 20300 2488
rect 19517 2483 19583 2486
rect 20294 2484 20300 2486
rect 20364 2484 20370 2548
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 20300 27236 20364 27300
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20300 22264 20364 22268
rect 20300 22208 20350 22264
rect 20350 22208 20364 22264
rect 20300 22204 20364 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 21588 20632 21652 20636
rect 21588 20576 21638 20632
rect 21638 20576 21652 20632
rect 21588 20572 21652 20576
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 20300 18668 20364 18732
rect 21036 18532 21100 18596
rect 21956 18532 22020 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 23244 17988 23308 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 21036 16764 21100 16828
rect 19380 16628 19444 16692
rect 20484 16492 20548 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 20116 16084 20180 16148
rect 21588 16084 21652 16148
rect 20852 15948 20916 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 20116 15676 20180 15740
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 19196 14860 19260 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 21956 14588 22020 14652
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 21036 13832 21100 13836
rect 21036 13776 21050 13832
rect 21050 13776 21100 13832
rect 21036 13772 21100 13776
rect 19196 13696 19260 13700
rect 19196 13640 19210 13696
rect 19210 13640 19260 13696
rect 19196 13636 19260 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 20300 13500 20364 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 14780 12820 14844 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 20484 11460 20548 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 26740 11188 26804 11252
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 20668 10780 20732 10844
rect 19196 10704 19260 10708
rect 19196 10648 19246 10704
rect 19246 10648 19260 10704
rect 19196 10644 19260 10648
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 20116 9964 20180 10028
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 17540 9616 17604 9620
rect 17540 9560 17554 9616
rect 17554 9560 17604 9616
rect 17540 9556 17604 9560
rect 20116 9420 20180 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 17540 8740 17604 8804
rect 20852 8740 20916 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 19196 8468 19260 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 25820 7516 25884 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 21036 6836 21100 6900
rect 28028 6836 28092 6900
rect 23244 6700 23308 6764
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 26740 6156 26804 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 14780 3980 14844 4044
rect 20116 3980 20180 4044
rect 20300 4040 20364 4044
rect 20300 3984 20350 4040
rect 20350 3984 20364 4040
rect 20300 3980 20364 3984
rect 28028 3980 28092 4044
rect 25820 3844 25884 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19380 3300 19444 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 20668 2892 20732 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 20300 2484 20364 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 20299 27300 20365 27301
rect 20299 27236 20300 27300
rect 20364 27236 20365 27300
rect 20299 27235 20365 27236
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 20302 22269 20362 27235
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 20299 22268 20365 22269
rect 20299 22204 20300 22268
rect 20364 22204 20365 22268
rect 20299 22203 20365 22204
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 21587 20636 21653 20637
rect 21587 20572 21588 20636
rect 21652 20572 21653 20636
rect 21587 20571 21653 20572
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20299 18732 20365 18733
rect 20299 18668 20300 18732
rect 20364 18668 20365 18732
rect 20299 18667 20365 18668
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19379 16692 19445 16693
rect 19379 16628 19380 16692
rect 19444 16628 19445 16692
rect 19379 16627 19445 16628
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 19195 14924 19261 14925
rect 19195 14860 19196 14924
rect 19260 14860 19261 14924
rect 19195 14859 19261 14860
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 19198 13701 19258 14859
rect 19195 13700 19261 13701
rect 19195 13636 19196 13700
rect 19260 13636 19261 13700
rect 19195 13635 19261 13636
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 14779 12884 14845 12885
rect 14779 12820 14780 12884
rect 14844 12820 14845 12884
rect 14779 12819 14845 12820
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 14782 4045 14842 12819
rect 19195 10708 19261 10709
rect 19195 10644 19196 10708
rect 19260 10644 19261 10708
rect 19195 10643 19261 10644
rect 17539 9620 17605 9621
rect 17539 9556 17540 9620
rect 17604 9556 17605 9620
rect 17539 9555 17605 9556
rect 17542 8805 17602 9555
rect 17539 8804 17605 8805
rect 17539 8740 17540 8804
rect 17604 8740 17605 8804
rect 17539 8739 17605 8740
rect 19198 8533 19258 10643
rect 19195 8532 19261 8533
rect 19195 8468 19196 8532
rect 19260 8468 19261 8532
rect 19195 8467 19261 8468
rect 14779 4044 14845 4045
rect 14779 3980 14780 4044
rect 14844 3980 14845 4044
rect 14779 3979 14845 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 19382 3365 19442 16627
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 20115 16148 20181 16149
rect 20115 16084 20116 16148
rect 20180 16084 20181 16148
rect 20115 16083 20181 16084
rect 20118 15741 20178 16083
rect 20115 15740 20181 15741
rect 20115 15676 20116 15740
rect 20180 15676 20181 15740
rect 20115 15675 20181 15676
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 20118 10029 20178 15675
rect 20302 13565 20362 18667
rect 21035 18596 21101 18597
rect 21035 18532 21036 18596
rect 21100 18532 21101 18596
rect 21035 18531 21101 18532
rect 21038 16829 21098 18531
rect 21035 16828 21101 16829
rect 21035 16764 21036 16828
rect 21100 16764 21101 16828
rect 21035 16763 21101 16764
rect 20483 16556 20549 16557
rect 20483 16492 20484 16556
rect 20548 16492 20549 16556
rect 20483 16491 20549 16492
rect 20299 13564 20365 13565
rect 20299 13500 20300 13564
rect 20364 13500 20365 13564
rect 20299 13499 20365 13500
rect 20486 11525 20546 16491
rect 21590 16149 21650 20571
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 21955 18596 22021 18597
rect 21955 18532 21956 18596
rect 22020 18532 22021 18596
rect 21955 18531 22021 18532
rect 21587 16148 21653 16149
rect 21587 16084 21588 16148
rect 21652 16084 21653 16148
rect 21587 16083 21653 16084
rect 20851 16012 20917 16013
rect 20851 15948 20852 16012
rect 20916 15948 20917 16012
rect 20851 15947 20917 15948
rect 20483 11524 20549 11525
rect 20483 11460 20484 11524
rect 20548 11460 20549 11524
rect 20483 11459 20549 11460
rect 20667 10844 20733 10845
rect 20667 10780 20668 10844
rect 20732 10780 20733 10844
rect 20667 10779 20733 10780
rect 20115 10028 20181 10029
rect 20115 9964 20116 10028
rect 20180 9964 20181 10028
rect 20115 9963 20181 9964
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 20115 9484 20181 9485
rect 20115 9420 20116 9484
rect 20180 9420 20181 9484
rect 20115 9419 20181 9420
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 3364 19445 3365
rect 19379 3300 19380 3364
rect 19444 3300 19445 3364
rect 19379 3299 19445 3300
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 20118 4045 20178 9419
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 20299 4044 20365 4045
rect 20299 3980 20300 4044
rect 20364 3980 20365 4044
rect 20299 3979 20365 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 20302 2549 20362 3979
rect 20670 2957 20730 10779
rect 20854 8805 20914 15947
rect 21958 14653 22018 18531
rect 23243 18052 23309 18053
rect 23243 17988 23244 18052
rect 23308 17988 23309 18052
rect 23243 17987 23309 17988
rect 21955 14652 22021 14653
rect 21955 14588 21956 14652
rect 22020 14588 22021 14652
rect 21955 14587 22021 14588
rect 21035 13836 21101 13837
rect 21035 13772 21036 13836
rect 21100 13772 21101 13836
rect 21035 13771 21101 13772
rect 20851 8804 20917 8805
rect 20851 8740 20852 8804
rect 20916 8740 20917 8804
rect 20851 8739 20917 8740
rect 21038 6901 21098 13771
rect 21035 6900 21101 6901
rect 21035 6836 21036 6900
rect 21100 6836 21101 6900
rect 21035 6835 21101 6836
rect 23246 6765 23306 17987
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 26739 11252 26805 11253
rect 26739 11188 26740 11252
rect 26804 11188 26805 11252
rect 26739 11187 26805 11188
rect 25819 7580 25885 7581
rect 25819 7516 25820 7580
rect 25884 7516 25885 7580
rect 25819 7515 25885 7516
rect 23243 6764 23309 6765
rect 23243 6700 23244 6764
rect 23308 6700 23309 6764
rect 23243 6699 23309 6700
rect 25822 3909 25882 7515
rect 26742 6221 26802 11187
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 28027 6900 28093 6901
rect 28027 6836 28028 6900
rect 28092 6836 28093 6900
rect 28027 6835 28093 6836
rect 26739 6220 26805 6221
rect 26739 6156 26740 6220
rect 26804 6156 26805 6220
rect 26739 6155 26805 6156
rect 28030 4045 28090 6835
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 28027 4044 28093 4045
rect 28027 3980 28028 4044
rect 28092 3980 28093 4044
rect 28027 3979 28093 3980
rect 25819 3908 25885 3909
rect 25819 3844 25820 3908
rect 25884 3844 25885 3908
rect 25819 3843 25885 3844
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20667 2956 20733 2957
rect 20667 2892 20668 2956
rect 20732 2892 20733 2956
rect 20667 2891 20733 2892
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 20299 2548 20365 2549
rect 20299 2484 20300 2548
rect 20364 2484 20365 2548
rect 20299 2483 20365 2484
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 26404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 17480 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1644511149
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1644511149
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1644511149
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1644511149
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1644511149
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_206
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1644511149
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1644511149
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_341
timestamp 1644511149
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1644511149
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1644511149
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1644511149
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1644511149
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1644511149
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_285
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_314
timestamp 1644511149
transform 1 0 29992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1644511149
transform 1 0 30728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1644511149
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1644511149
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_371
timestamp 1644511149
transform 1 0 35236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1644511149
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_157
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_268
timestamp 1644511149
transform 1 0 25760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_278
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp 1644511149
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1644511149
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_319
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_341
timestamp 1644511149
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_351
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1644511149
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1644511149
transform 1 0 37720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1644511149
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1644511149
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_126
timestamp 1644511149
transform 1 0 12696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1644511149
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_265
timestamp 1644511149
transform 1 0 25484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_286
timestamp 1644511149
transform 1 0 27416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1644511149
transform 1 0 29624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_343
timestamp 1644511149
transform 1 0 32660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_351
timestamp 1644511149
transform 1 0 33396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1644511149
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_377
timestamp 1644511149
transform 1 0 35788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_383
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_397
timestamp 1644511149
transform 1 0 37628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_35
timestamp 1644511149
transform 1 0 4324 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1644511149
transform 1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_52
timestamp 1644511149
transform 1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1644511149
transform 1 0 6624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_106
timestamp 1644511149
transform 1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1644511149
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1644511149
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1644511149
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_256
timestamp 1644511149
transform 1 0 24656 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_268
timestamp 1644511149
transform 1 0 25760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1644511149
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1644511149
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_291
timestamp 1644511149
transform 1 0 27876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1644511149
transform 1 0 30084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_319
timestamp 1644511149
transform 1 0 30452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_326
timestamp 1644511149
transform 1 0 31096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1644511149
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_339
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_352
timestamp 1644511149
transform 1 0 33488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1644511149
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_370
timestamp 1644511149
transform 1 0 35144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_379
timestamp 1644511149
transform 1 0 35972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_383
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_397
timestamp 1644511149
transform 1 0 37628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1644511149
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1644511149
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1644511149
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_79
timestamp 1644511149
transform 1 0 8372 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1644511149
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_118
timestamp 1644511149
transform 1 0 11960 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_140
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1644511149
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1644511149
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1644511149
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1644511149
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_206
timestamp 1644511149
transform 1 0 20056 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_212
timestamp 1644511149
transform 1 0 20608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1644511149
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1644511149
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_238
timestamp 1644511149
transform 1 0 23000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_246
timestamp 1644511149
transform 1 0 23736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_253
timestamp 1644511149
transform 1 0 24380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_260
timestamp 1644511149
transform 1 0 25024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_267
timestamp 1644511149
transform 1 0 25668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1644511149
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_284
timestamp 1644511149
transform 1 0 27232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_292
timestamp 1644511149
transform 1 0 27968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_298
timestamp 1644511149
transform 1 0 28520 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_304
timestamp 1644511149
transform 1 0 29072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1644511149
transform 1 0 29624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_319
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_326
timestamp 1644511149
transform 1 0 31096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1644511149
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_342
timestamp 1644511149
transform 1 0 32568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_351
timestamp 1644511149
transform 1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_358
timestamp 1644511149
transform 1 0 34040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_365
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1644511149
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_398
timestamp 1644511149
transform 1 0 37720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1644511149
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1644511149
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1644511149
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1644511149
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1644511149
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_123
timestamp 1644511149
transform 1 0 12420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1644511149
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_147
timestamp 1644511149
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1644511149
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_161
timestamp 1644511149
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_168
timestamp 1644511149
transform 1 0 16560 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_174
timestamp 1644511149
transform 1 0 17112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1644511149
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_218
timestamp 1644511149
transform 1 0 21160 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1644511149
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_293
timestamp 1644511149
transform 1 0 28060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_297
timestamp 1644511149
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_316
timestamp 1644511149
transform 1 0 30176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_329
timestamp 1644511149
transform 1 0 31372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_340
timestamp 1644511149
transform 1 0 32384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_349
timestamp 1644511149
transform 1 0 33212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1644511149
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_373
timestamp 1644511149
transform 1 0 35420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_380
timestamp 1644511149
transform 1 0 36064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1644511149
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_394
timestamp 1644511149
transform 1 0 37352 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_398
timestamp 1644511149
transform 1 0 37720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1644511149
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1644511149
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_67
timestamp 1644511149
transform 1 0 7268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1644511149
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1644511149
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1644511149
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_143
timestamp 1644511149
transform 1 0 14260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_157
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1644511149
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_180
timestamp 1644511149
transform 1 0 17664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1644511149
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_247
timestamp 1644511149
transform 1 0 23828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp 1644511149
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_260
timestamp 1644511149
transform 1 0 25024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_269
timestamp 1644511149
transform 1 0 25852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_297
timestamp 1644511149
transform 1 0 28428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1644511149
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_325
timestamp 1644511149
transform 1 0 31004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_345
timestamp 1644511149
transform 1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_360
timestamp 1644511149
transform 1 0 34224 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_368
timestamp 1644511149
transform 1 0 34960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1644511149
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_396
timestamp 1644511149
transform 1 0 37536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1644511149
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1644511149
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_35
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_42
timestamp 1644511149
transform 1 0 4968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1644511149
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1644511149
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_94
timestamp 1644511149
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1644511149
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_110
timestamp 1644511149
transform 1 0 11224 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp 1644511149
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1644511149
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1644511149
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_167
timestamp 1644511149
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_171
timestamp 1644511149
transform 1 0 16836 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_205
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_211
timestamp 1644511149
transform 1 0 20516 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_216
timestamp 1644511149
transform 1 0 20976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1644511149
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_234
timestamp 1644511149
transform 1 0 22632 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1644511149
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_270
timestamp 1644511149
transform 1 0 25944 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1644511149
transform 1 0 26496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_283
timestamp 1644511149
transform 1 0 27140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_293
timestamp 1644511149
transform 1 0 28060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_325
timestamp 1644511149
transform 1 0 31004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_351
timestamp 1644511149
transform 1 0 33396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1644511149
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_381
timestamp 1644511149
transform 1 0 36156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_391
timestamp 1644511149
transform 1 0 37076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1644511149
transform 1 0 37720 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1644511149
transform 1 0 38456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_6
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1644511149
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1644511149
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1644511149
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1644511149
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1644511149
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_92
timestamp 1644511149
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_118
timestamp 1644511149
transform 1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_140
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_146
timestamp 1644511149
transform 1 0 14536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1644511149
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_186
timestamp 1644511149
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1644511149
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_232
timestamp 1644511149
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 1644511149
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_240
timestamp 1644511149
transform 1 0 23184 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_250
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_268
timestamp 1644511149
transform 1 0 25760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_272
timestamp 1644511149
transform 1 0 26128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_294
timestamp 1644511149
transform 1 0 28152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_301
timestamp 1644511149
transform 1 0 28796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_321
timestamp 1644511149
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_330
timestamp 1644511149
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_353
timestamp 1644511149
transform 1 0 33580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1644511149
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_396
timestamp 1644511149
transform 1 0 37536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1644511149
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1644511149
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1644511149
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1644511149
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_59
timestamp 1644511149
transform 1 0 6532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1644511149
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1644511149
transform 1 0 14352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1644511149
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_175
timestamp 1644511149
transform 1 0 17204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_186
timestamp 1644511149
transform 1 0 18216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1644511149
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_212
timestamp 1644511149
transform 1 0 20608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1644511149
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1644511149
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_269
timestamp 1644511149
transform 1 0 25852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_275
timestamp 1644511149
transform 1 0 26404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_283
timestamp 1644511149
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1644511149
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_335
timestamp 1644511149
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_342
timestamp 1644511149
transform 1 0 32568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_349
timestamp 1644511149
transform 1 0 33212 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1644511149
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_371
timestamp 1644511149
transform 1 0 35236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_378
timestamp 1644511149
transform 1 0 35880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_385
timestamp 1644511149
transform 1 0 36524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_393
timestamp 1644511149
transform 1 0 37260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_402
timestamp 1644511149
transform 1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1644511149
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_8
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1644511149
transform 1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1644511149
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 1644511149
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1644511149
transform 1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1644511149
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1644511149
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1644511149
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1644511149
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1644511149
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_124
timestamp 1644511149
transform 1 0 12512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1644511149
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1644511149
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1644511149
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1644511149
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_228
timestamp 1644511149
transform 1 0 22080 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_234
timestamp 1644511149
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1644511149
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1644511149
transform 1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_268
timestamp 1644511149
transform 1 0 25760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1644511149
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1644511149
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_328
timestamp 1644511149
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_340
timestamp 1644511149
transform 1 0 32384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_351
timestamp 1644511149
transform 1 0 33396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_358
timestamp 1644511149
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_365
timestamp 1644511149
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_372 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_16
timestamp 1644511149
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_48
timestamp 1644511149
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1644511149
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1644511149
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_90
timestamp 1644511149
transform 1 0 9384 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_96
timestamp 1644511149
transform 1 0 9936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1644511149
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1644511149
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_159
timestamp 1644511149
transform 1 0 15732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1644511149
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_216
timestamp 1644511149
transform 1 0 20976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_234
timestamp 1644511149
transform 1 0 22632 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_242
timestamp 1644511149
transform 1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_270
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_278
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_286
timestamp 1644511149
transform 1 0 27416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1644511149
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1644511149
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_312
timestamp 1644511149
transform 1 0 29808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_319
timestamp 1644511149
transform 1 0 30452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_326
timestamp 1644511149
transform 1 0 31096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_340
timestamp 1644511149
transform 1 0 32384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_347
timestamp 1644511149
transform 1 0 33028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_354
timestamp 1644511149
transform 1 0 33672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1644511149
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_65
timestamp 1644511149
transform 1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1644511149
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1644511149
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1644511149
transform 1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1644511149
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1644511149
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1644511149
transform 1 0 18768 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_200
timestamp 1644511149
transform 1 0 19504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_231
timestamp 1644511149
transform 1 0 22356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1644511149
transform 1 0 23184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1644511149
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_258
timestamp 1644511149
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_267
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_288
timestamp 1644511149
transform 1 0 27600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_295
timestamp 1644511149
transform 1 0 28244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_315
timestamp 1644511149
transform 1 0 30084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_322
timestamp 1644511149
transform 1 0 30728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1644511149
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_347
timestamp 1644511149
transform 1 0 33028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_354
timestamp 1644511149
transform 1 0 33672 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_366
timestamp 1644511149
transform 1 0 34776 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_378
timestamp 1644511149
transform 1 0 35880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1644511149
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1644511149
transform 1 0 6440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1644511149
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1644511149
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1644511149
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_104
timestamp 1644511149
transform 1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1644511149
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1644511149
transform 1 0 11960 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp 1644511149
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1644511149
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_146
timestamp 1644511149
transform 1 0 14536 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1644511149
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1644511149
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_180
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_186
timestamp 1644511149
transform 1 0 18216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1644511149
transform 1 0 20056 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_214
timestamp 1644511149
transform 1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_274
timestamp 1644511149
transform 1 0 26312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1644511149
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_297
timestamp 1644511149
transform 1 0 28428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_312
timestamp 1644511149
transform 1 0 29808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_319
timestamp 1644511149
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_326
timestamp 1644511149
transform 1 0 31096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1644511149
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_70
timestamp 1644511149
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1644511149
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1644511149
transform 1 0 8740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1644511149
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_122
timestamp 1644511149
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1644511149
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_142
timestamp 1644511149
transform 1 0 14168 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1644511149
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_182
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1644511149
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_206
timestamp 1644511149
transform 1 0 20056 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1644511149
transform 1 0 20700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_228
timestamp 1644511149
transform 1 0 22080 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_232
timestamp 1644511149
transform 1 0 22448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_238
timestamp 1644511149
transform 1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_250
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1644511149
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_285
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_313
timestamp 1644511149
transform 1 0 29900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_318
timestamp 1644511149
transform 1 0 30360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1644511149
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_88
timestamp 1644511149
transform 1 0 9200 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1644511149
transform 1 0 11224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1644511149
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1644511149
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_213
timestamp 1644511149
transform 1 0 20700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_228
timestamp 1644511149
transform 1 0 22080 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_234
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1644511149
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_258
timestamp 1644511149
transform 1 0 24840 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_272
timestamp 1644511149
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_284
timestamp 1644511149
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1644511149
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1644511149
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_312
timestamp 1644511149
transform 1 0 29808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_319
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1644511149
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1644511149
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_118
timestamp 1644511149
transform 1 0 11960 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1644511149
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1644511149
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1644511149
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_202
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1644511149
transform 1 0 20516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_238
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_264
timestamp 1644511149
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_284
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_314
timestamp 1644511149
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 1644511149
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1644511149
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_88
timestamp 1644511149
transform 1 0 9200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_96
timestamp 1644511149
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1644511149
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_107
timestamp 1644511149
transform 1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_115
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1644511149
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_126
timestamp 1644511149
transform 1 0 12696 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1644511149
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_157
timestamp 1644511149
transform 1 0 15548 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_214
timestamp 1644511149
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1644511149
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_257
timestamp 1644511149
transform 1 0 24748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_266
timestamp 1644511149
transform 1 0 25576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_280
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_312
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_324
timestamp 1644511149
transform 1 0 30912 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_336
timestamp 1644511149
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_348
timestamp 1644511149
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1644511149
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1644511149
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_212
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_216
timestamp 1644511149
transform 1 0 20976 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_234
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1644511149
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_289
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_315
timestamp 1644511149
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp 1644511149
transform 1 0 31188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1644511149
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_116
timestamp 1644511149
transform 1 0 11776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_120
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1644511149
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1644511149
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1644511149
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_151
timestamp 1644511149
transform 1 0 14996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_176
timestamp 1644511149
transform 1 0 17296 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1644511149
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_226
timestamp 1644511149
transform 1 0 21896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1644511149
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1644511149
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1644511149
transform 1 0 11960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1644511149
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_134
timestamp 1644511149
transform 1 0 13432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1644511149
transform 1 0 15456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1644511149
transform 1 0 17204 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_183
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_262
timestamp 1644511149
transform 1 0 25208 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1644511149
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1644511149
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1644511149
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_116
timestamp 1644511149
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_127
timestamp 1644511149
transform 1 0 12788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1644511149
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_270
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_296
timestamp 1644511149
transform 1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1644511149
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_337
timestamp 1644511149
transform 1 0 32108 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_349
timestamp 1644511149
transform 1 0 33212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1644511149
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1644511149
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1644511149
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1644511149
transform 1 0 13524 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_143
timestamp 1644511149
transform 1 0 14260 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1644511149
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1644511149
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_228
timestamp 1644511149
transform 1 0 22080 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_246
timestamp 1644511149
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1644511149
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1644511149
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_298
timestamp 1644511149
transform 1 0 28520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_322
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1644511149
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1644511149
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_116
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_156
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_171
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_187
timestamp 1644511149
transform 1 0 18308 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_227
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_298
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1644511149
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1644511149
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_102
timestamp 1644511149
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1644511149
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1644511149
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1644511149
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_138
timestamp 1644511149
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_144
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_197
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_230
timestamp 1644511149
transform 1 0 22264 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_246
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_266
timestamp 1644511149
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1644511149
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_285
timestamp 1644511149
transform 1 0 27324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_297
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_304
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_310
timestamp 1644511149
transform 1 0 29624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_318
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_344
timestamp 1644511149
transform 1 0 32752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_352
timestamp 1644511149
transform 1 0 33488 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_364
timestamp 1644511149
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_376
timestamp 1644511149
transform 1 0 35696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1644511149
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1644511149
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp 1644511149
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1644511149
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_206
timestamp 1644511149
transform 1 0 20056 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1644511149
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_227
timestamp 1644511149
transform 1 0 21988 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_235
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1644511149
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1644511149
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_319
timestamp 1644511149
transform 1 0 30452 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_325
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_348
timestamp 1644511149
transform 1 0 33120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1644511149
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1644511149
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_127
timestamp 1644511149
transform 1 0 12788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_135
timestamp 1644511149
transform 1 0 13524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1644511149
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1644511149
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_263
timestamp 1644511149
transform 1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1644511149
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_284
timestamp 1644511149
transform 1 0 27232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_292
timestamp 1644511149
transform 1 0 27968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1644511149
transform 1 0 32660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1644511149
transform 1 0 33764 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1644511149
transform 1 0 34868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1644511149
transform 1 0 35972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_108
timestamp 1644511149
transform 1 0 11040 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_128
timestamp 1644511149
transform 1 0 12880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_152
timestamp 1644511149
transform 1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_219
timestamp 1644511149
transform 1 0 21252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1644511149
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1644511149
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1644511149
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_299
timestamp 1644511149
transform 1 0 28612 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_328
timestamp 1644511149
transform 1 0 31280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_334
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1644511149
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_129
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_153
timestamp 1644511149
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1644511149
transform 1 0 22816 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1644511149
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_257
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_265
timestamp 1644511149
transform 1 0 25484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_271
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_288
timestamp 1644511149
transform 1 0 27600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1644511149
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_343
timestamp 1644511149
transform 1 0 32660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_351
timestamp 1644511149
transform 1 0 33396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_128
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1644511149
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1644511149
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_231
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_328
timestamp 1644511149
transform 1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1644511149
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_122
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_178
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_191
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1644511149
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1644511149
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_300
timestamp 1644511149
transform 1 0 28704 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_304
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_311
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_319
timestamp 1644511149
transform 1 0 30452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_350
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_357
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_369
timestamp 1644511149
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_381
timestamp 1644511149
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1644511149
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_210
timestamp 1644511149
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_241
timestamp 1644511149
transform 1 0 23276 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_262
timestamp 1644511149
transform 1 0 25208 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_283
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_290
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_316
timestamp 1644511149
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_336
timestamp 1644511149
transform 1 0 32016 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_349
timestamp 1644511149
transform 1 0 33212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1644511149
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_373
timestamp 1644511149
transform 1 0 35420 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_385
timestamp 1644511149
transform 1 0 36524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_397
timestamp 1644511149
transform 1 0 37628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1644511149
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_130
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_152
timestamp 1644511149
transform 1 0 15088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_207
timestamp 1644511149
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_230
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_238
timestamp 1644511149
transform 1 0 23000 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_255
timestamp 1644511149
transform 1 0 24564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_269
timestamp 1644511149
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_288
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_296
timestamp 1644511149
transform 1 0 28336 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_322
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_368
timestamp 1644511149
transform 1 0 34960 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_380
timestamp 1644511149
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_129
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1644511149
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_147
timestamp 1644511149
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1644511149
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_159
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_167
timestamp 1644511149
transform 1 0 16468 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1644511149
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_215
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_223
timestamp 1644511149
transform 1 0 21620 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1644511149
transform 1 0 21988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1644511149
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_286
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1644511149
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_344
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_353
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_175
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_183
timestamp 1644511149
transform 1 0 17940 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_200
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_208
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_230
timestamp 1644511149
transform 1 0 22264 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1644511149
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_250
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1644511149
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_298
timestamp 1644511149
transform 1 0 28520 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_310
timestamp 1644511149
transform 1 0 29624 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_320
timestamp 1644511149
transform 1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1644511149
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_343
timestamp 1644511149
transform 1 0 32660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_351
timestamp 1644511149
transform 1 0 33396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_368
timestamp 1644511149
transform 1 0 34960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_376
timestamp 1644511149
transform 1 0 35696 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_117
timestamp 1644511149
transform 1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1644511149
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_156
timestamp 1644511149
transform 1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1644511149
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_222
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_257
timestamp 1644511149
transform 1 0 24748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_279
timestamp 1644511149
transform 1 0 26772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_334
timestamp 1644511149
transform 1 0 31832 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_349
timestamp 1644511149
transform 1 0 33212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1644511149
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_141
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1644511149
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_191
timestamp 1644511149
transform 1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_197
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1644511149
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_248
timestamp 1644511149
transform 1 0 23920 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_252
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_303
timestamp 1644511149
transform 1 0 28980 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_344
timestamp 1644511149
transform 1 0 32752 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_366
timestamp 1644511149
transform 1 0 34776 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_378
timestamp 1644511149
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1644511149
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 1644511149
transform 1 0 11776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_125
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_176
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_202
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_215
timestamp 1644511149
transform 1 0 20884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_290
timestamp 1644511149
transform 1 0 27784 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_296
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1644511149
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_322
timestamp 1644511149
transform 1 0 30728 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_330
timestamp 1644511149
transform 1 0 31464 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_336
timestamp 1644511149
transform 1 0 32016 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_346
timestamp 1644511149
transform 1 0 32936 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_368
timestamp 1644511149
transform 1 0 34960 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_380
timestamp 1644511149
transform 1 0 36064 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_392
timestamp 1644511149
transform 1 0 37168 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_404
timestamp 1644511149
transform 1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_132
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_138
timestamp 1644511149
transform 1 0 13800 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_148
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_178
timestamp 1644511149
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1644511149
transform 1 0 23460 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1644511149
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_299
timestamp 1644511149
transform 1 0 28612 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_307
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_315
timestamp 1644511149
transform 1 0 30084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_346
timestamp 1644511149
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_358
timestamp 1644511149
transform 1 0 34040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_365
timestamp 1644511149
transform 1 0 34684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_377
timestamp 1644511149
transform 1 0 35788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1644511149
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_125
timestamp 1644511149
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1644511149
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1644511149
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_200
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_207
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_216
timestamp 1644511149
transform 1 0 20976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_234
timestamp 1644511149
transform 1 0 22632 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_238
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_260
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_276
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_284
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_331
timestamp 1644511149
transform 1 0 31556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_150
timestamp 1644511149
transform 1 0 14904 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_192
timestamp 1644511149
transform 1 0 18768 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_235
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_244
timestamp 1644511149
transform 1 0 23552 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_248
timestamp 1644511149
transform 1 0 23920 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_253
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_265
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_284
timestamp 1644511149
transform 1 0 27232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_292
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_320
timestamp 1644511149
transform 1 0 30544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1644511149
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_345
timestamp 1644511149
transform 1 0 32844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_357
timestamp 1644511149
transform 1 0 33948 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_369
timestamp 1644511149
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1644511149
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_117
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_123
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_157
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_208
timestamp 1644511149
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_262
timestamp 1644511149
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_282
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_328
timestamp 1644511149
transform 1 0 31280 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_348
timestamp 1644511149
transform 1 0 33120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_136
timestamp 1644511149
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_174
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_187
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_207
timestamp 1644511149
transform 1 0 20148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_211
timestamp 1644511149
transform 1 0 20516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_228
timestamp 1644511149
transform 1 0 22080 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_232
timestamp 1644511149
transform 1 0 22448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_246
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_268
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_301
timestamp 1644511149
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_313
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_325
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1644511149
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_150
timestamp 1644511149
transform 1 0 14904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_168
timestamp 1644511149
transform 1 0 16560 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_172
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_231
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_239
timestamp 1644511149
transform 1 0 23092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_257
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_295
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1644511149
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1644511149
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_182
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_206
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_213
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_238
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_260
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1644511149
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_309
timestamp 1644511149
transform 1 0 29532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_321
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1644511149
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_171
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1644511149
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_219
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_227
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_256
timestamp 1644511149
transform 1 0 24656 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_174
timestamp 1644511149
transform 1 0 17112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_189
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1644511149
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_250
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_176
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_204
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1644511149
transform 1 0 21896 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1644511149
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_157
timestamp 1644511149
transform 1 0 15548 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_172
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1644511149
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1644511149
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_228
timestamp 1644511149
transform 1 0 22080 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_240
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_252
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_264
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_175
timestamp 1644511149
transform 1 0 17204 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1644511149
transform 1 0 18032 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 1644511149
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1644511149
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_217
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1644511149
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_200
timestamp 1644511149
transform 1 0 19504 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_212
timestamp 1644511149
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_224
timestamp 1644511149
transform 1 0 21712 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_236
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_201
timestamp 1644511149
transform 1 0 19596 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_206
timestamp 1644511149
transform 1 0 20056 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_218
timestamp 1644511149
transform 1 0 21160 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_47
timestamp 1644511149
transform 1 0 5428 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1644511149
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1644511149
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_155
timestamp 1644511149
transform 1 0 15364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1644511149
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_264
timestamp 1644511149
transform 1 0 25392 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1644511149
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1644511149
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_373
timestamp 1644511149
transform 1 0 35420 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_385
timestamp 1644511149
transform 1 0 36524 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_391
timestamp 1644511149
transform 1 0 37076 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0782_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0783_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5336 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0784_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0785_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0786_
timestamp 1644511149
transform 1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0787_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9108 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0788_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0789_
timestamp 1644511149
transform 1 0 10672 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1644511149
transform 1 0 12052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0791_
timestamp 1644511149
transform 1 0 14996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0792_
timestamp 1644511149
transform 1 0 13616 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0793_
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_2  _0794_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0795_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0796_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0797_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0798_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0799_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0800_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1644511149
transform 1 0 23552 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0803_
timestamp 1644511149
transform 1 0 33304 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0804_
timestamp 1644511149
transform 1 0 30728 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0805_
timestamp 1644511149
transform 1 0 31372 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0806_
timestamp 1644511149
transform 1 0 31096 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_2  _0807_
timestamp 1644511149
transform 1 0 32384 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1644511149
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0809_
timestamp 1644511149
transform 1 0 31096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _0810_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0811_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32752 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0812_
timestamp 1644511149
transform 1 0 33488 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0813_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0814_
timestamp 1644511149
transform 1 0 32200 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0815_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33212 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _0816_
timestamp 1644511149
transform 1 0 33764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _0817_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0818_
timestamp 1644511149
transform 1 0 30912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0819_
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0820_
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_1  _0821_
timestamp 1644511149
transform 1 0 31096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0822_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0823_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0824_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29992 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0825_
timestamp 1644511149
transform 1 0 30084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0826_
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0827_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0828_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0829_
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1644511149
transform 1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0832_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0834_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31832 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0835_
timestamp 1644511149
transform 1 0 32752 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0836_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0837_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _0838_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _0839_
timestamp 1644511149
transform 1 0 27140 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0840_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0841_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0842_
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0843_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0845_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0846_
timestamp 1644511149
transform 1 0 35052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0848_
timestamp 1644511149
transform 1 0 25944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0849_
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0850_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0851_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _0852_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0853_
timestamp 1644511149
transform 1 0 26128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0854_
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0855_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0856_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0857_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21712 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0858_
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0860_
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0862_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _0863_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0864_
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0865_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0867_
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0868_
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0869_
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0870_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0871_
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0873_
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0874_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0876_
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0877_
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0878_
timestamp 1644511149
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0879_
timestamp 1644511149
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0880_
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 1644511149
transform 1 0 19780 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0882_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0883_
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp 1644511149
transform 1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0888_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0889_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0891_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0893_
timestamp 1644511149
transform 1 0 6532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0894_
timestamp 1644511149
transform 1 0 14444 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0895_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0896_
timestamp 1644511149
transform 1 0 21068 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0899_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0900_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0901_
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0902_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0903_
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0904_
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1644511149
transform 1 0 22080 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0906_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1644511149
transform 1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1644511149
transform 1 0 24472 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1644511149
transform 1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1644511149
transform 1 0 23552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0911_
timestamp 1644511149
transform 1 0 24564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0912_
timestamp 1644511149
transform 1 0 23000 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0915_
timestamp 1644511149
transform 1 0 22448 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0916_
timestamp 1644511149
transform 1 0 22632 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 1644511149
transform 1 0 22724 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 1644511149
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1644511149
transform 1 0 23552 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0922_
timestamp 1644511149
transform 1 0 25576 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0924_
timestamp 1644511149
transform 1 0 25116 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0925_
timestamp 1644511149
transform 1 0 25392 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0928_
timestamp 1644511149
transform 1 0 26680 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0929_
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 1644511149
transform 1 0 26036 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0931_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1644511149
transform 1 0 24932 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0935_
timestamp 1644511149
transform 1 0 23368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1644511149
transform 1 0 23460 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1644511149
transform 1 0 24104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1644511149
transform 1 0 24748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 1644511149
transform 1 0 26496 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0940_
timestamp 1644511149
transform 1 0 26680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1644511149
transform 1 0 24932 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1644511149
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0943_
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0945_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0946_
timestamp 1644511149
transform 1 0 24472 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1644511149
transform 1 0 24196 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1644511149
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0949_
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0950_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0951_
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0952_
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1644511149
transform 1 0 26128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0955_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _0956_
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0958_
timestamp 1644511149
transform 1 0 26128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0960_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0963_
timestamp 1644511149
transform 1 0 27508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0964_
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0967_
timestamp 1644511149
transform 1 0 26128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 1644511149
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _0970_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0972_
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0974_
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0975_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1644511149
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0977_
timestamp 1644511149
transform 1 0 24104 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0978_
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0979_
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0981_
timestamp 1644511149
transform 1 0 25760 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0982_
timestamp 1644511149
transform 1 0 26496 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1644511149
transform 1 0 26772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1644511149
transform 1 0 30544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0985_
timestamp 1644511149
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1644511149
transform 1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0989_
timestamp 1644511149
transform 1 0 29532 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1644511149
transform 1 0 33856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0991_
timestamp 1644511149
transform 1 0 28612 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1644511149
transform 1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0993_
timestamp 1644511149
transform 1 0 29992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1644511149
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1644511149
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0997_
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1644511149
transform 1 0 31464 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform 1 0 32292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1001_
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1644511149
transform 1 0 32936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1003_
timestamp 1644511149
transform 1 0 32384 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1644511149
transform 1 0 36432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1005_
timestamp 1644511149
transform 1 0 32752 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1644511149
transform 1 0 37076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1644511149
transform 1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1644511149
transform 1 0 33120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1009_
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1011_
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 37904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1013_
timestamp 1644511149
transform 1 0 35328 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1015_
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 1644511149
transform 1 0 35788 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1644511149
transform 1 0 36984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1644511149
transform 1 0 33304 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1020_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1644511149
transform 1 0 37904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1644511149
transform 1 0 37812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1024_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1026_
timestamp 1644511149
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1027_
timestamp 1644511149
transform 1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1029_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1030_
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1644511149
transform 1 0 13340 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1644511149
transform 1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1033_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1644511149
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1035_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1644511149
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1038_
timestamp 1644511149
transform 1 0 15364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1039_
timestamp 1644511149
transform 1 0 12880 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1644511149
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1041_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1644511149
transform 1 0 10212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1043_
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1048_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1644511149
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1644511149
transform 1 0 12328 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1644511149
transform 1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1054_
timestamp 1644511149
transform 1 0 10580 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1644511149
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1644511149
transform 1 0 29716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1059_
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1060_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1061_
timestamp 1644511149
transform 1 0 16008 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1644511149
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1063_
timestamp 1644511149
transform 1 0 17664 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkinv_2  _1064_
timestamp 1644511149
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1065_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1066_
timestamp 1644511149
transform 1 0 23000 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1067_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1068_
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1069_
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1072_
timestamp 1644511149
transform 1 0 24932 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1073_
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1644511149
transform 1 0 22632 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1075_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1076_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1077_
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1078_
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1079_
timestamp 1644511149
transform 1 0 15272 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1080_
timestamp 1644511149
transform 1 0 15272 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1081_
timestamp 1644511149
transform 1 0 16008 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1082_
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1083_
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1084_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1086_
timestamp 1644511149
transform 1 0 20976 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1644511149
transform 1 0 15272 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1089_
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1090_
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1644511149
transform 1 0 18216 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1093_
timestamp 1644511149
transform 1 0 12144 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1644511149
transform 1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1095_
timestamp 1644511149
transform 1 0 17204 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1096_
timestamp 1644511149
transform 1 0 16744 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1098_
timestamp 1644511149
transform 1 0 17020 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1644511149
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1101_
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1102_
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1104_
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1107_
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1108_
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1111_
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1112_
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1644511149
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1644511149
transform 1 0 14904 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1116_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1117_
timestamp 1644511149
transform 1 0 14720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1118_
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1644511149
transform 1 0 17296 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1644511149
transform 1 0 9016 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1123_
timestamp 1644511149
transform 1 0 18124 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1124_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1644511149
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1644511149
transform 1 0 8096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1127_
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1644511149
transform 1 0 19780 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1130_
timestamp 1644511149
transform 1 0 12420 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1131_
timestamp 1644511149
transform 1 0 18124 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1644511149
transform 1 0 17756 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1644511149
transform 1 0 17572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1134_
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1644511149
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1137_
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1140_
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1644511149
transform 1 0 18124 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1142_
timestamp 1644511149
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1143_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1644511149
transform 1 0 18584 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1644511149
transform 1 0 19320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1146_
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1147_
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1148_
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1644511149
transform 1 0 3864 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1150_
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1151_
timestamp 1644511149
transform 1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1644511149
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1154_
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1155_
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1158_
timestamp 1644511149
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1159_
timestamp 1644511149
transform 1 0 6440 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1160_
timestamp 1644511149
transform 1 0 7084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1162_
timestamp 1644511149
transform 1 0 8464 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1163_
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1644511149
transform 1 0 4784 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1165_
timestamp 1644511149
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1166_
timestamp 1644511149
transform 1 0 9384 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1167_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1168_
timestamp 1644511149
transform 1 0 5612 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1644511149
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1170_
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1171_
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1173_
timestamp 1644511149
transform 1 0 5888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1644511149
transform 1 0 5060 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1176_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1182_
timestamp 1644511149
transform 1 0 10120 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1183_
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1184_
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 1644511149
transform 1 0 7820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1188_
timestamp 1644511149
transform 1 0 7728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1190_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1191_
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1644511149
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1194_
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1195_
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1196_
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1644511149
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1198_
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1199_
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1203_
timestamp 1644511149
transform 1 0 9568 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1204_
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1206_
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1644511149
transform 1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1209_
timestamp 1644511149
transform 1 0 10948 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1212_
timestamp 1644511149
transform 1 0 9936 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1644511149
transform 1 0 10580 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1218_
timestamp 1644511149
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1219_
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1220_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1644511149
transform 1 0 12788 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1223_
timestamp 1644511149
transform 1 0 11316 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1224_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1226_
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1227_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1228_
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1229_
timestamp 1644511149
transform 1 0 14720 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1230_
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1231_
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1234_
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1644511149
transform 1 0 12788 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1644511149
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1237_
timestamp 1644511149
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1238_
timestamp 1644511149
transform 1 0 12972 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1240_
timestamp 1644511149
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1241_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1644511149
transform 1 0 12880 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1243_
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1244_
timestamp 1644511149
transform 1 0 12972 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1245_
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1247_
timestamp 1644511149
transform 1 0 14260 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1250_
timestamp 1644511149
transform 1 0 14628 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 14444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1253_
timestamp 1644511149
transform 1 0 14904 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1644511149
transform 1 0 16376 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1256_
timestamp 1644511149
transform 1 0 14904 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1644511149
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1259_
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1260_
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1262_
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1264_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1265_
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1266_
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1267_
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1269_
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1270_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _1271_
timestamp 1644511149
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1272_
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1273_
timestamp 1644511149
transform 1 0 25392 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1274_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1275_
timestamp 1644511149
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1276_
timestamp 1644511149
transform 1 0 29808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1277_
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1278_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1279_
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1280_
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1644511149
transform 1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1282_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1283_
timestamp 1644511149
transform 1 0 27600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1644511149
transform 1 0 27048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1286_
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1287_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1644511149
transform 1 0 28520 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1644511149
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _1290_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1291_
timestamp 1644511149
transform 1 0 27048 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1292_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1293_
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1295_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1296_
timestamp 1644511149
transform 1 0 31096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1644511149
transform 1 0 30912 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1299_
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1301_
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1302_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1303_
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1304_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1306_
timestamp 1644511149
transform 1 0 30544 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1307_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1308_
timestamp 1644511149
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1309_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1310_
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1311_
timestamp 1644511149
transform 1 0 33672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1312_
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1313_
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1314_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1315_
timestamp 1644511149
transform 1 0 32384 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1316_
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1317_
timestamp 1644511149
transform 1 0 32476 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1644511149
transform 1 0 35328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1321_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1644511149
transform 1 0 33764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1323_
timestamp 1644511149
transform 1 0 32292 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1324_
timestamp 1644511149
transform 1 0 32568 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1325_
timestamp 1644511149
transform 1 0 32200 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1326_
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1328_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1644511149
transform 1 0 33304 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1332_
timestamp 1644511149
transform 1 0 19412 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1333_
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1334_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1335_
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1336_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1337_
timestamp 1644511149
transform 1 0 16836 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1338_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1339_
timestamp 1644511149
transform 1 0 13248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1340_
timestamp 1644511149
transform 1 0 16560 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1342_
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1343_
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1344_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1345_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1346_
timestamp 1644511149
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1347_
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1348_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1349_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1350_
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1351_
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1352_
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1353_
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1354_
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1355_
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1356_
timestamp 1644511149
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1357_
timestamp 1644511149
transform 1 0 13616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1358_
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1359_
timestamp 1644511149
transform 1 0 14628 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1360_
timestamp 1644511149
transform 1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1361_
timestamp 1644511149
transform 1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1362_
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1644511149
transform 1 0 16836 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1364_
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1365_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1366_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1367_
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1368_
timestamp 1644511149
transform 1 0 17940 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1369_
timestamp 1644511149
transform 1 0 18216 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1370_
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1371_
timestamp 1644511149
transform 1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1372_
timestamp 1644511149
transform 1 0 18032 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1373_
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1374_
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1375_
timestamp 1644511149
transform 1 0 20056 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1376_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1377_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1378_
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1379_
timestamp 1644511149
transform 1 0 16744 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1380_
timestamp 1644511149
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1381_
timestamp 1644511149
transform 1 0 20884 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1644511149
transform 1 0 20240 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1383_
timestamp 1644511149
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1384_
timestamp 1644511149
transform 1 0 26772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1385_
timestamp 1644511149
transform 1 0 21988 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1386_
timestamp 1644511149
transform 1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1387_
timestamp 1644511149
transform 1 0 26036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1388_
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1390_
timestamp 1644511149
transform 1 0 27784 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1644511149
transform 1 0 28980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1392_
timestamp 1644511149
transform 1 0 22724 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1644511149
transform 1 0 20424 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1644511149
transform 1 0 27600 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1397_
timestamp 1644511149
transform 1 0 30084 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1398_
timestamp 1644511149
transform 1 0 25392 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1644511149
transform 1 0 30176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1644511149
transform 1 0 28612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1644511149
transform 1 0 28060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1402_
timestamp 1644511149
transform 1 0 28428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1403_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1644511149
transform 1 0 27968 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1644511149
transform 1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1406_
timestamp 1644511149
transform 1 0 30452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1644511149
transform 1 0 27600 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1644511149
transform 1 0 28428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp 1644511149
transform 1 0 31464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1410_
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1411_
timestamp 1644511149
transform 1 0 30176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1412_
timestamp 1644511149
transform 1 0 24656 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1644511149
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1414_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1415_
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1416_
timestamp 1644511149
transform 1 0 29256 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1417_
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1418_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1419_
timestamp 1644511149
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1420_
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1421_
timestamp 1644511149
transform 1 0 29716 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1644511149
transform 1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1423_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 1644511149
transform 1 0 31004 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1425_
timestamp 1644511149
transform 1 0 32108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1426_
timestamp 1644511149
transform 1 0 30544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1644511149
transform 1 0 34408 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1428_
timestamp 1644511149
transform 1 0 31464 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1429_
timestamp 1644511149
transform 1 0 32384 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1430_
timestamp 1644511149
transform 1 0 32752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1431_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1432_
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 33396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1434_
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1435_
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1644511149
transform 1 0 35052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1437_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1438_
timestamp 1644511149
transform 1 0 35512 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1440_
timestamp 1644511149
transform 1 0 36524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1441_
timestamp 1644511149
transform 1 0 34960 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1442_
timestamp 1644511149
transform 1 0 36248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1443_
timestamp 1644511149
transform 1 0 35788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1445_
timestamp 1644511149
transform 1 0 24472 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1446_
timestamp 1644511149
transform 1 0 24564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1447_
timestamp 1644511149
transform 1 0 21712 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1448_
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1451_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1452_
timestamp 1644511149
transform 1 0 22080 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1453_
timestamp 1644511149
transform 1 0 25944 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1454_
timestamp 1644511149
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1455_
timestamp 1644511149
transform 1 0 24748 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1456_
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1457_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1458_
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1460_
timestamp 1644511149
transform 1 0 28704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1462_
timestamp 1644511149
transform 1 0 29624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1463_
timestamp 1644511149
transform 1 0 27784 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1464_
timestamp 1644511149
transform 1 0 25300 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1465_
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1466_
timestamp 1644511149
transform 1 0 23276 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1467_
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1468_
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1469_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1470_
timestamp 1644511149
transform 1 0 26220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1471_
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1472_
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1473_
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1474_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1475_
timestamp 1644511149
transform 1 0 25208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1476_
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1477_
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1478_
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1479_
timestamp 1644511149
transform 1 0 25208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1480_
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1481_
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1482_
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1483_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1484_
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1485_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1486_
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 1644511149
transform 1 0 22908 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1489_
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1490_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1491_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1492_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1493_
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1644511149
transform 1 0 15272 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1495_
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 1644511149
transform 1 0 15824 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1497_
timestamp 1644511149
transform 1 0 15272 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1498_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1499_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1501_
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1502_
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1503_
timestamp 1644511149
transform 1 0 18308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1644511149
transform 1 0 16468 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1506_
timestamp 1644511149
transform 1 0 15640 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1508_
timestamp 1644511149
transform 1 0 20608 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1509_
timestamp 1644511149
transform 1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1510_
timestamp 1644511149
transform 1 0 16928 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1511_
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1512_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1513_
timestamp 1644511149
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1515_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1516_
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1644511149
transform 1 0 17848 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 1644511149
transform 1 0 16744 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1644511149
transform 1 0 18308 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1520_
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1521_
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1522_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1644511149
transform 1 0 14076 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1524_
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1525_
timestamp 1644511149
transform 1 0 15272 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 1644511149
transform 1 0 13984 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1527_
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1528_
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1529_
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1530_
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1532_
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1644511149
transform 1 0 14260 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1534_
timestamp 1644511149
transform 1 0 16100 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1535_
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1536_
timestamp 1644511149
transform 1 0 15916 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1537_
timestamp 1644511149
transform 1 0 20608 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1538_
timestamp 1644511149
transform 1 0 19872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 1644511149
transform 1 0 12788 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1540_
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1541_
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1644511149
transform 1 0 12144 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1543_
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1544_
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1545_
timestamp 1644511149
transform 1 0 13892 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1546_
timestamp 1644511149
transform 1 0 12972 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1547_
timestamp 1644511149
transform 1 0 12144 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1549_
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1550_
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1644511149
transform 1 0 14444 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1552_
timestamp 1644511149
transform 1 0 12972 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1554_
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1555_
timestamp 1644511149
transform 1 0 19320 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1556_
timestamp 1644511149
transform 1 0 18400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1644511149
transform 1 0 12972 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1559_
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1560_
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1561_
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1644511149
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1563_
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1644511149
transform 1 0 17664 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1644511149
transform 1 0 17940 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1566_
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1567_
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1568_
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1570_
timestamp 1644511149
transform 1 0 19320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform 1 0 19780 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1575_
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1644511149
transform 1 0 17848 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1644511149
transform 1 0 17572 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1580_
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1583_
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1586_
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1588_
timestamp 1644511149
transform 1 0 22264 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1589_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1590_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1592_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1593_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1595_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1596_
timestamp 1644511149
transform 1 0 24564 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1599_
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1600_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1644511149
transform 1 0 9476 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1644511149
transform 1 0 12052 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1644511149
transform 1 0 9476 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1644511149
transform 1 0 9476 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1644511149
transform 1 0 9476 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1644511149
transform 1 0 11408 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1644511149
transform 1 0 11592 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1644511149
transform 1 0 22356 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1612_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1644511149
transform 1 0 24104 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1644511149
transform 1 0 16192 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1615_
timestamp 1644511149
transform 1 0 16928 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1617_
timestamp 1644511149
transform 1 0 18032 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1618_
timestamp 1644511149
transform 1 0 14536 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1619_
timestamp 1644511149
transform 1 0 19596 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1644511149
transform 1 0 12696 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1621_
timestamp 1644511149
transform 1 0 20884 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1644511149
transform 1 0 13432 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1644511149
transform 1 0 15824 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1644511149
transform 1 0 19872 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1644511149
transform 1 0 17020 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1644511149
transform 1 0 6532 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1634_
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1644511149
transform 1 0 4232 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1644511149
transform 1 0 4324 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1644511149
transform 1 0 4140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1644511149
transform 1 0 4048 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1644511149
transform 1 0 5520 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1644511149
transform 1 0 6900 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1644511149
transform 1 0 8004 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1644511149
transform 1 0 9384 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1644511149
transform 1 0 9016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1644511149
transform 1 0 9752 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1644511149
transform 1 0 9844 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1644511149
transform 1 0 11592 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1644511149
transform 1 0 10948 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1644511149
transform 1 0 11684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1644511149
transform 1 0 12512 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1644511149
transform 1 0 14260 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1644511149
transform 1 0 14536 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1663_
timestamp 1644511149
transform 1 0 22264 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1644511149
transform 1 0 27416 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1644511149
transform 1 0 29072 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1644511149
transform 1 0 29808 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1644511149
transform 1 0 31648 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1644511149
transform 1 0 33304 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1644511149
transform 1 0 32108 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1644511149
transform 1 0 15640 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1644511149
transform 1 0 14352 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1644511149
transform 1 0 14260 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1685_
timestamp 1644511149
transform 1 0 18124 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1687_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 21160 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 22080 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 24840 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 28612 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 22448 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1644511149
transform 1 0 28520 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 24472 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 27140 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1644511149
transform 1 0 28612 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1644511149
transform 1 0 26220 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1644511149
transform 1 0 27600 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 27508 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 24472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 29992 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 31924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1644511149
transform 1 0 33488 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1644511149
transform 1 0 33948 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1644511149
transform 1 0 35236 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1644511149
transform 1 0 35144 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1727_
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1644511149
transform 1 0 29256 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1644511149
transform 1 0 22540 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1644511149
transform 1 0 22724 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1644511149
transform 1 0 25576 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1644511149
transform 1 0 17204 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1644511149
transform 1 0 14628 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1644511149
transform 1 0 12144 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1644511149
transform 1 0 12788 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1644511149
transform 1 0 15824 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1644511149
transform 1 0 20424 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1644511149
transform 1 0 17112 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1644511149
transform 1 0 19872 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1758__90 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1759__91
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_CLK
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_CLK
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_CLK
timestamp 1644511149
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_CLK
timestamp 1644511149
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_CLK
timestamp 1644511149
transform 1 0 28612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_CLK
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_CLK
timestamp 1644511149
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_CLK
timestamp 1644511149
transform 1 0 12880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_CLK
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_CLK
timestamp 1644511149
transform 1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_CLK
timestamp 1644511149
transform 1 0 26036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_CLK
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_CLK
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_CLK
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_CLK
timestamp 1644511149
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_CLK
timestamp 1644511149
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_CLK
timestamp 1644511149
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_CLK
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_CLK
timestamp 1644511149
transform 1 0 11224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_CLK
timestamp 1644511149
transform 1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_CLK
timestamp 1644511149
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_CLK
timestamp 1644511149
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_CLK
timestamp 1644511149
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_CLK
timestamp 1644511149
transform 1 0 24472 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_CLK
timestamp 1644511149
transform 1 0 33764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_CLK
timestamp 1644511149
transform 1 0 29992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_CLK
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_CLK
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_CLK
timestamp 1644511149
transform 1 0 28336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_CLK
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 15364 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 30176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 30728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 31464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 32752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 31464 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 22080 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 33396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1644511149
transform 1 0 5060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1644511149
transform 1 0 28244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 33948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 37352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 25024 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 35052 0 1 46784
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 570 0 626 800 6 RST_N
port 1 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 slave_ack_o
port 2 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 slave_adr_i[0]
port 3 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 slave_adr_i[10]
port 4 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 slave_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 slave_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 slave_adr_i[13]
port 7 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 slave_adr_i[14]
port 8 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 slave_adr_i[15]
port 9 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 slave_adr_i[16]
port 10 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 slave_adr_i[17]
port 11 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 slave_adr_i[18]
port 12 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 slave_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 slave_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 slave_adr_i[20]
port 15 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 slave_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 slave_adr_i[22]
port 17 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 slave_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 slave_adr_i[24]
port 19 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 slave_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 slave_adr_i[26]
port 21 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 slave_adr_i[27]
port 22 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 slave_adr_i[28]
port 23 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 slave_adr_i[29]
port 24 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 slave_adr_i[2]
port 25 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 slave_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 slave_adr_i[31]
port 27 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 slave_adr_i[3]
port 28 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 slave_adr_i[4]
port 29 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 slave_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 slave_adr_i[6]
port 31 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 slave_adr_i[7]
port 32 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 slave_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 slave_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 938 0 994 800 6 slave_cyc_i
port 35 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 slave_dat_i[0]
port 36 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 slave_dat_i[10]
port 37 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 slave_dat_i[11]
port 38 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 slave_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 slave_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 slave_dat_i[14]
port 41 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 slave_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 slave_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 slave_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 slave_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 slave_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 slave_dat_i[1]
port 47 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 slave_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 slave_dat_i[21]
port 49 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 slave_dat_i[22]
port 50 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 slave_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 slave_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 slave_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 slave_dat_i[26]
port 54 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 slave_dat_i[27]
port 55 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 slave_dat_i[28]
port 56 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 slave_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 slave_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 slave_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 slave_dat_i[31]
port 60 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 slave_dat_i[3]
port 61 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 slave_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 slave_dat_i[5]
port 63 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 slave_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 slave_dat_i[7]
port 65 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 slave_dat_i[8]
port 66 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 slave_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 slave_dat_o[0]
port 68 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 slave_dat_o[10]
port 69 nsew signal tristate
rlabel metal2 s 24582 0 24638 800 6 slave_dat_o[11]
port 70 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 slave_dat_o[12]
port 71 nsew signal tristate
rlabel metal2 s 26054 0 26110 800 6 slave_dat_o[13]
port 72 nsew signal tristate
rlabel metal2 s 26882 0 26938 800 6 slave_dat_o[14]
port 73 nsew signal tristate
rlabel metal2 s 27618 0 27674 800 6 slave_dat_o[15]
port 74 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 slave_dat_o[16]
port 75 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 slave_dat_o[17]
port 76 nsew signal tristate
rlabel metal2 s 29826 0 29882 800 6 slave_dat_o[18]
port 77 nsew signal tristate
rlabel metal2 s 30562 0 30618 800 6 slave_dat_o[19]
port 78 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 slave_dat_o[1]
port 79 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 slave_dat_o[20]
port 80 nsew signal tristate
rlabel metal2 s 32034 0 32090 800 6 slave_dat_o[21]
port 81 nsew signal tristate
rlabel metal2 s 32770 0 32826 800 6 slave_dat_o[22]
port 82 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 slave_dat_o[23]
port 83 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 slave_dat_o[24]
port 84 nsew signal tristate
rlabel metal2 s 34978 0 35034 800 6 slave_dat_o[25]
port 85 nsew signal tristate
rlabel metal2 s 35714 0 35770 800 6 slave_dat_o[26]
port 86 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 slave_dat_o[27]
port 87 nsew signal tristate
rlabel metal2 s 37186 0 37242 800 6 slave_dat_o[28]
port 88 nsew signal tristate
rlabel metal2 s 37922 0 37978 800 6 slave_dat_o[29]
port 89 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 slave_dat_o[2]
port 90 nsew signal tristate
rlabel metal2 s 38658 0 38714 800 6 slave_dat_o[30]
port 91 nsew signal tristate
rlabel metal2 s 39394 0 39450 800 6 slave_dat_o[31]
port 92 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 slave_dat_o[3]
port 93 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 slave_dat_o[4]
port 94 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 slave_dat_o[5]
port 95 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 slave_dat_o[6]
port 96 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 slave_dat_o[7]
port 97 nsew signal tristate
rlabel metal2 s 22374 0 22430 800 6 slave_dat_o[8]
port 98 nsew signal tristate
rlabel metal2 s 23110 0 23166 800 6 slave_dat_o[9]
port 99 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 slave_err_o
port 100 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 slave_rty_o
port 101 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 slave_sel_i[0]
port 102 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 slave_sel_i[1]
port 103 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 slave_sel_i[2]
port 104 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 slave_sel_i[3]
port 105 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 slave_stb_i
port 106 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 slave_we_i
port 107 nsew signal input
rlabel metal2 s 4986 49200 5042 50000 6 spiMaster_miso
port 108 nsew signal input
rlabel metal2 s 14922 49200 14978 50000 6 spiMaster_mosi
port 109 nsew signal tristate
rlabel metal2 s 24950 49200 25006 50000 6 spiMaster_mosi_oe
port 110 nsew signal tristate
rlabel metal2 s 34978 49200 35034 50000 6 spiMaster_sclk
port 111 nsew signal tristate
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 112 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 112 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 113 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
